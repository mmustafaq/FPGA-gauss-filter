library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.pcg.all;


entity sdram is

port(

CLOCK_50: IN STD_LOGIC;
SW: IN STD_LOGIC_VECTOR(9 downto 0);
----------------VGA-Interface---------------------
VGA_B,VGA_G,VGA_R : OUT STD_LOGIC_VECTOR(7 downto 0);
VGA_CLK,VGA_BLANK_N,VGA_HS,VGA_VS,VGA_SYNC_N: OUT STD_LOGIC;
LEDR: OUT STD_LOGIC_VECTOR(9 downto 0);
KEY: IN STD_LOGIC_VECTOR(3 downto 0);
------------------SDRAM---------------------------
DRAM_ADDR: OUT STD_LOGIC_VECTOR(12 downto 0);
DRAM_BA: OUT STD_LOGIC_VECTOR(1 downto 0);
DRAM_CAS_N: OUT STD_LOGIC;
DRAM_CKE: OUT STD_LOGIC;
DRAM_CLK: OUT STD_LOGIC;
DRAM_CS_N: OUT STD_LOGIC;
DRAM_DQ: INOUT STD_LOGIC_VECTOR(15 downto 0);
DRAM_RAS_N: OUT STD_LOGIC;
DRAM_WE_N: OUT STD_LOGIC;
DRAM_LDQM,DRAM_UDQM: OUT STD_LOGIC
);


end sdram;


architecture  main of sdram is
TYPE STAGES IS (ST0,ST1);
SIGNAL BUFF_CTRL: STAGES:=ST0;
---------------------------test signals----------------------------
type Array4096 is array (0 to 65535) of integer;
constant ROM: Array4096 :=(
153,153,153,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,155,154,155,154,154,154,155,155,154,155,155,155,154,155,155,154,154,154,155,154,155,155,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,154,155,155,154,155,154,155,155,155,154,155,155,155,155,155,155,155,155,155,156,156,156,156,156,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,158,158,157,158,157,157,158,158,158,156,151,153,153,154,155,155,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,158,158,158,158,158,157,158,158,158,158,159,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,159,160,160,160,159,160,161,160,160,161,160,160,161,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,160,160,161,161,160,160,160,160,160,159,157,160,121,157,163,159,164,152,101,116,165,155,100,
154,154,154,154,154,155,154,154,155,155,154,155,155,155,155,155,155,156,156,155,156,156,155,155,155,156,155,155,155,155,155,156,156,156,156,155,155,155,155,155,155,156,155,155,155,156,156,156,156,155,155,155,154,154,155,155,155,155,155,156,155,156,156,155,155,156,156,155,155,156,156,156,156,156,156,156,156,157,156,157,157,157,157,157,156,156,157,157,157,157,157,158,157,157,158,157,157,158,158,158,157,158,158,158,157,158,158,158,158,158,159,158,158,159,158,158,158,158,158,157,157,158,155,155,156,155,156,157,157,157,157,157,158,158,158,158,158,158,158,158,158,159,159,158,159,158,159,158,158,158,158,158,158,159,158,159,159,159,159,159,159,159,159,159,159,160,159,159,160,160,160,160,160,160,160,160,160,160,160,160,161,161,160,161,161,161,160,161,160,161,161,161,161,161,160,161,161,161,161,161,161,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,160,161,161,161,161,161,160,160,160,161,160,161,161,161,160,163,159,153,161,154,153,161,134,149,160,124,152,121,
154,155,155,155,155,155,155,155,156,155,156,156,156,156,156,156,156,156,156,156,156,156,156,156,155,155,155,155,156,156,156,156,157,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,155,155,155,155,154,155,156,156,157,157,156,156,157,156,156,156,156,156,156,156,156,157,157,156,157,156,157,157,157,157,157,158,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,158,158,158,158,158,158,159,158,159,159,160,159,159,158,159,159,159,160,159,157,157,156,157,157,157,157,158,157,157,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,159,159,159,159,159,159,159,159,159,160,159,159,159,160,160,160,159,160,160,160,160,161,161,160,161,161,160,160,161,162,161,161,161,161,161,162,162,162,161,161,162,162,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,163,162,171,156,134,159,159,191,184,200,128,158,164,150,
156,155,155,155,156,156,156,156,156,156,156,157,157,157,157,157,156,156,157,157,157,157,157,156,157,157,156,156,156,157,157,156,157,157,156,157,157,157,157,157,157,157,157,157,156,157,156,157,157,156,157,156,156,156,157,156,155,155,157,157,157,157,156,157,157,157,156,157,156,157,157,157,157,157,158,158,157,157,157,157,157,158,157,157,158,158,157,158,158,158,159,159,158,158,159,159,159,159,159,159,159,159,159,159,159,159,158,159,159,159,159,159,159,159,159,159,160,159,159,159,160,159,159,158,158,157,158,157,157,158,157,159,158,159,159,159,159,159,159,159,159,160,160,160,160,159,160,160,160,160,160,159,160,159,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,160,161,161,161,161,162,161,162,162,162,162,162,162,162,162,162,161,162,162,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,161,162,162,162,161,162,162,161,162,162,166,158,170,167,158,163,170,168,147,165,161,152,175,143,
156,156,156,155,156,156,157,157,157,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,156,157,157,157,158,157,157,157,157,157,158,157,157,157,158,158,157,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,159,160,160,160,160,160,160,160,159,159,159,159,158,158,158,158,159,159,159,159,159,159,160,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,160,160,161,161,161,161,160,160,161,161,162,163,162,161,161,162,161,162,161,162,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,162,162,162,162,162,162,162,162,162,162,163,163,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,162,162,164,167,162,162,162,162,162,162,162,163,162,162,163,162,162,162,163,162,163,164,164,149,139,123,164,172,163,160,185,169,106,112,160,134,109,
156,156,156,156,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,157,157,157,158,158,157,157,158,157,158,158,158,158,158,157,157,158,158,158,158,158,158,158,158,157,158,158,157,157,158,157,157,158,158,158,157,158,157,158,158,157,158,158,158,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,159,160,160,160,160,160,160,160,160,160,160,160,161,160,160,160,160,160,160,160,160,160,159,159,159,159,159,159,160,160,160,160,159,160,160,160,161,160,160,160,160,161,161,161,160,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,161,162,162,161,162,162,162,162,162,162,162,162,162,162,163,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,162,164,163,163,163,159,177,155,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,157,163,133,66,101,194,180,163,163,181,109,57,152,129,134,172,
157,157,156,157,158,157,157,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,158,157,158,158,158,158,158,158,158,158,158,158,159,158,158,158,158,159,158,158,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,158,159,159,159,159,158,159,159,159,158,159,159,159,159,159,159,159,159,159,159,160,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,161,161,161,161,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,160,160,160,161,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,161,162,162,162,161,162,162,162,162,162,162,163,162,162,162,162,162,163,163,163,162,163,163,163,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,163,163,163,164,163,163,163,164,163,163,163,163,163,163,163,163,164,165,170,164,162,162,163,163,163,163,163,163,163,163,161,165,163,163,163,163,163,163,163,163,163,161,164,164,163,155,160,159,176,125,139,161,174,135,160,139,156,123,136,182,143,183,147,
157,158,158,158,158,158,158,158,159,158,158,158,158,158,158,158,158,159,158,159,159,159,159,159,159,159,159,158,159,158,159,159,158,158,158,158,159,159,159,159,158,158,159,159,159,159,159,158,158,158,158,158,159,159,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,159,159,159,159,159,160,160,160,160,160,159,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,161,161,161,162,162,162,162,161,161,162,161,162,162,161,161,161,161,161,161,160,161,161,161,161,161,161,161,161,161,161,161,162,163,162,162,162,162,162,162,162,162,162,162,162,162,162,163,162,163,162,162,163,163,163,163,163,163,162,162,163,163,163,163,164,163,163,163,163,163,163,163,163,164,164,163,164,164,164,164,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,150,165,161,169,164,164,164,164,164,164,162,164,164,157,165,165,164,164,164,164,164,164,174,164,164,165,163,154,164,125,165,95,184,164,167,166,183,175,200,156,103,142,109,172,144,
158,158,158,159,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,159,159,159,159,159,159,159,160,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,159,159,159,159,159,159,159,160,160,159,160,160,160,160,160,160,160,160,160,160,159,160,160,160,161,160,160,161,161,161,161,161,161,162,162,161,161,161,162,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,161,161,161,161,161,161,161,161,162,162,161,161,162,163,164,163,163,164,164,163,163,163,163,163,163,163,163,164,163,163,163,164,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,164,164,164,164,164,164,164,165,165,165,165,165,165,162,164,165,170,162,166,165,165,165,169,161,173,162,164,165,166,165,166,165,165,163,168,168,157,165,164,165,165,164,164,134,161,169,132,175,170,175,154,127,181,153,159,124,102,90,129,
158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,159,160,159,159,159,160,160,159,160,159,159,159,159,159,160,160,160,159,159,160,160,160,159,159,160,159,159,159,159,159,159,160,159,159,160,160,159,160,159,159,160,160,160,160,160,160,160,160,160,160,160,160,161,161,160,160,160,160,160,160,160,161,160,161,160,161,160,161,161,161,161,161,161,162,161,162,162,162,162,162,161,162,162,162,162,162,162,162,162,162,163,164,163,163,163,163,163,162,162,162,162,163,163,163,163,163,162,162,162,163,162,162,163,162,162,162,162,162,163,162,163,163,164,164,164,164,164,164,164,164,164,164,164,163,164,164,164,163,164,164,164,164,165,164,164,164,164,165,165,164,164,164,164,164,164,164,164,164,165,165,164,164,165,164,164,164,164,165,164,165,165,164,164,165,165,165,164,165,165,165,165,165,165,165,165,164,165,165,164,165,166,165,185,162,150,168,161,168,158,167,165,166,165,163,163,165,165,166,167,167,166,166,167,166,158,152,165,165,165,166,165,166,161,157,167,190,143,127,177,181,119,179,120,126,102,62,143,163,
159,159,159,159,159,159,159,159,159,160,159,159,160,159,160,160,160,160,160,160,160,160,160,161,160,160,160,160,160,160,160,160,160,160,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,160,160,160,160,161,161,161,160,161,161,160,161,161,160,161,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,161,162,162,162,162,162,163,162,163,162,162,163,163,163,164,163,164,164,164,163,164,164,164,163,163,164,164,164,163,163,164,163,165,164,164,163,163,163,163,162,163,163,164,163,163,163,163,163,163,164,165,164,164,165,165,165,165,165,165,164,164,165,165,165,165,164,164,165,164,164,164,165,165,165,163,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,166,166,166,166,165,166,165,165,166,165,165,165,166,165,165,166,166,165,165,166,166,166,115,143,179,170,165,159,176,163,167,164,165,166,164,164,166,169,167,167,96,166,166,153,170,137,162,166,166,166,166,166,160,174,149,145,171,174,190,89,153,176,154,140,131,105,120,134,113,
160,159,159,160,160,160,161,161,160,161,160,160,160,161,160,160,160,160,160,160,160,160,160,161,161,161,161,161,160,161,161,161,160,160,161,160,160,161,162,160,160,160,160,160,161,161,161,161,161,161,160,161,161,161,161,161,161,161,161,160,160,161,161,161,161,161,161,161,161,161,161,160,161,161,161,161,161,161,161,161,161,161,162,161,162,162,162,162,162,162,162,163,162,163,163,163,163,164,162,164,162,163,164,164,164,164,164,164,164,164,164,164,165,165,165,164,164,165,165,164,164,164,164,164,164,165,164,164,165,165,164,164,164,164,165,165,164,164,164,165,164,165,165,165,165,165,165,165,165,165,165,165,164,165,165,165,165,164,165,165,164,165,164,165,165,165,165,164,165,165,165,165,164,165,165,165,165,165,165,166,165,165,166,165,165,162,166,166,166,166,166,166,167,166,166,166,165,166,166,165,166,166,167,166,166,166,166,167,165,166,172,144,169,157,168,146,170,155,169,168,166,163,165,178,158,180,158,142,169,168,167,119,171,165,166,166,167,166,168,187,132,191,170,168,156,178,141,173,124,174,135,134,145,110,78,141,
160,160,160,160,161,160,161,161,161,162,161,161,161,161,162,161,161,161,161,161,161,161,161,161,162,162,161,161,162,162,162,162,162,161,162,162,161,161,161,161,161,161,162,162,161,161,161,161,161,162,161,161,161,162,161,162,162,161,162,162,162,162,162,162,162,163,162,162,162,162,161,162,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,163,162,162,164,163,164,164,165,164,164,164,165,165,164,165,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,165,165,165,165,165,165,165,165,166,164,165,165,166,166,165,166,166,165,165,165,165,165,165,166,165,166,165,165,165,165,165,165,165,166,165,166,166,165,165,165,166,166,166,166,166,165,166,165,165,165,165,165,166,166,167,167,167,166,166,166,166,166,166,166,167,167,167,167,167,167,166,167,167,167,167,167,167,167,167,167,168,166,167,167,173,167,140,205,115,142,134,156,169,172,170,169,167,169,176,171,161,164,156,128,164,167,166,168,167,167,165,167,172,166,131,138,142,161,191,174,159,156,165,195,130,119,103,184,142,161,
161,161,162,161,162,161,161,161,161,162,162,161,161,162,162,161,161,162,162,161,162,161,162,161,162,162,162,163,163,163,163,162,163,162,163,162,163,161,162,162,162,162,163,161,162,161,161,162,160,162,163,163,162,163,163,162,163,163,163,163,163,163,162,163,163,162,163,164,163,163,162,163,162,163,162,162,163,163,163,163,163,163,163,162,163,163,163,164,163,164,165,164,164,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,165,166,167,165,165,165,166,166,166,165,166,166,165,165,165,166,165,165,165,166,166,165,165,165,165,166,166,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,166,166,166,166,165,166,166,166,165,166,166,166,166,166,167,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,167,168,167,166,167,167,167,167,167,167,166,167,169,167,174,167,197,114,154,154,147,135,168,167,149,156,155,158,178,166,171,170,173,102,190,149,181,182,168,169,177,140,147,148,170,172,163,144,190,162,170,139,81,142,123,129,130,125,73,108,171,
161,162,162,162,162,162,163,163,162,162,162,163,163,163,162,163,163,163,163,163,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,162,162,162,163,163,162,163,163,163,163,163,163,163,163,163,164,164,164,164,163,163,164,163,164,163,163,164,163,162,163,163,164,163,163,164,164,163,163,164,164,164,164,164,164,164,165,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,166,166,166,166,166,166,166,167,167,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,166,167,167,167,167,167,166,166,167,167,167,167,167,167,166,167,167,167,167,167,167,166,166,166,166,166,167,167,168,168,167,168,167,167,168,167,167,167,168,168,168,168,168,168,168,168,168,168,167,167,167,167,167,161,169,166,162,171,167,167,140,152,150,146,171,125,177,175,89,186,116,172,149,170,130,142,167,166,175,134,122,169,179,158,173,129,158,143,150,157,174,123,147,177,132,183,178,183,194,145,103,191,163,110,
163,163,163,163,162,163,163,163,163,163,163,164,163,164,163,163,163,163,163,163,163,163,163,162,163,163,164,164,164,165,163,163,163,164,164,164,164,164,163,164,164,164,163,163,164,164,163,164,164,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,164,164,165,165,165,164,164,164,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,165,165,166,166,166,166,166,166,166,165,166,166,166,166,166,167,166,166,166,167,167,167,166,167,167,167,167,166,166,167,167,167,167,167,166,166,167,167,167,167,167,167,167,168,167,167,167,168,167,168,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,168,168,168,168,167,168,168,168,169,169,169,169,169,169,169,169,168,167,167,167,167,170,145,164,163,159,127,121,175,155,218,144,152,171,168,142,150,164,135,145,146,168,169,180,150,156,128,157,157,185,160,170,173,152,182,132,168,174,149,172,196,154,162,87,142,140,116,130,132,198,116,106,
163,163,163,163,163,164,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,163,165,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,164,165,165,165,165,165,165,165,165,165,165,165,165,165,164,165,165,165,165,165,165,165,165,165,165,165,166,165,165,166,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,167,168,167,167,167,167,166,168,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,167,167,168,168,168,167,167,167,167,167,167,168,167,168,168,168,168,169,168,168,169,169,168,169,169,169,169,169,169,169,169,170,169,169,169,169,167,167,167,165,170,166,161,178,97,132,170,167,163,151,152,144,160,180,103,136,86,81,130,107,125,161,169,93,168,128,149,121,75,164,183,177,181,180,182,174,159,186,169,118,133,163,154,124,239,89,127,125,167,153,
163,163,163,163,164,164,164,164,163,164,164,164,164,164,164,164,165,164,164,164,164,164,164,165,165,165,164,164,165,164,164,164,164,165,165,165,165,164,164,164,164,165,165,165,165,165,165,165,164,165,164,165,165,165,165,166,165,165,165,165,165,165,165,165,165,166,166,165,165,166,164,165,165,165,165,165,165,166,166,166,166,165,166,166,166,166,166,165,167,166,166,167,166,166,166,167,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,167,167,167,168,168,167,167,168,168,168,167,168,167,167,168,168,168,168,168,168,167,168,168,168,167,168,168,168,168,168,168,168,168,169,169,169,169,168,169,168,168,169,168,168,168,168,169,169,169,168,169,168,169,169,168,168,168,168,168,168,169,168,168,167,167,167,167,169,169,169,169,169,169,169,169,169,170,170,169,169,169,169,170,171,171,171,171,170,169,171,168,145,149,173,176,181,183,181,184,140,169,169,172,164,167,164,134,137,81,165,129,162,154,112,165,136,166,157,152,124,109,145,180,175,137,133,128,138,172,141,126,170,164,94,110,145,71,115,136,138,148,125,161,
164,164,164,163,164,164,165,165,165,164,164,164,164,164,165,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,165,165,165,165,165,165,165,165,165,166,165,165,165,165,165,165,166,166,166,166,165,166,166,166,166,165,166,166,165,165,166,166,165,166,166,166,165,165,166,166,166,166,166,166,166,166,166,166,167,166,167,166,167,166,167,167,167,167,167,167,167,167,167,168,168,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,168,168,168,169,168,168,168,168,170,168,168,169,168,169,169,169,169,168,168,168,169,169,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,169,169,169,169,169,169,169,170,169,169,169,169,169,169,168,168,170,170,169,169,169,169,170,170,170,170,170,170,170,168,172,171,170,171,170,171,171,171,171,177,171,174,179,158,149,167,168,180,160,186,154,217,110,189,190,139,179,110,142,187,119,127,98,119,165,165,165,146,125,187,80,113,152,118,128,178,172,196,170,149,133,134,116,75,107,93,137,179,115,98,133,123,
164,164,164,165,164,165,165,165,165,164,166,166,165,165,165,165,165,165,165,165,166,165,166,166,166,165,165,165,166,166,166,165,166,165,165,166,165,166,165,166,166,165,166,166,166,166,165,166,166,165,166,165,166,165,165,166,166,166,166,165,166,166,166,166,166,165,167,167,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,166,167,167,167,167,167,167,167,167,167,167,168,167,168,168,168,168,168,168,168,168,169,168,168,169,168,169,168,168,168,168,169,169,168,168,169,169,169,169,169,169,168,168,169,169,168,169,169,169,168,167,169,169,169,167,169,170,170,169,169,169,169,170,170,170,170,169,170,169,170,170,170,170,170,170,170,170,171,170,169,170,169,170,170,170,170,170,170,170,171,170,170,170,170,170,169,170,169,170,170,170,170,170,171,170,171,171,171,169,172,172,171,173,174,172,174,164,171,174,168,145,122,142,168,139,155,118,119,168,153,149,136,102,181,104,72,168,159,147,84,149,97,126,135,166,167,186,182,143,150,152,131,166,151,163,159,107,140,160,76,137,133,97,115,90,115,151,146,154,
165,165,165,165,165,165,165,165,166,165,166,166,166,166,166,166,166,166,166,166,165,166,166,166,165,166,166,166,165,165,166,166,166,166,166,166,166,166,166,166,166,165,166,166,166,166,166,166,166,166,166,166,166,166,167,166,166,166,166,166,166,167,166,166,167,166,167,167,167,167,166,166,166,167,167,167,167,167,166,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,168,169,169,168,170,169,170,170,169,169,170,169,169,169,169,170,169,169,170,170,169,170,170,170,170,171,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,170,170,170,171,171,171,170,171,170,171,170,171,170,171,171,171,171,171,171,171,171,171,171,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,174,172,173,176,172,172,171,176,151,125,180,151,165,188,152,153,134,165,176,100,151,185,186,167,119,92,137,182,140,138,134,154,151,177,145,160,126,145,115,141,132,105,145,163,146,142,145,114,148,184,87,166,95,133,142,124,130,154,167,106,
165,165,165,165,165,166,166,166,166,166,166,166,165,166,166,165,166,166,166,166,166,166,167,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,166,167,167,166,166,166,166,166,166,167,167,167,167,166,166,167,167,167,167,167,168,167,167,167,167,167,167,167,167,167,167,167,167,168,168,167,167,167,167,168,167,168,168,168,167,168,168,169,168,169,168,169,169,169,169,169,169,169,170,169,170,170,170,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,169,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,170,171,170,171,171,171,171,171,171,171,171,171,171,171,172,171,171,172,171,171,171,171,171,171,171,172,172,172,172,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,173,172,173,172,173,173,175,174,200,139,162,84,137,144,148,128,141,116,173,147,74,175,141,69,191,166,184,187,115,142,179,148,150,154,182,112,125,144,198,59,109,181,141,160,160,143,176,128,174,173,126,140,158,144,108,156,160,147,
166,166,166,165,165,165,166,166,166,166,166,166,166,167,166,166,167,167,167,167,167,167,167,167,167,167,166,167,167,167,167,167,166,166,166,167,166,167,167,167,167,167,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,168,169,169,169,169,169,170,170,170,170,170,170,171,170,170,171,170,170,171,171,171,171,171,170,170,170,170,170,170,171,171,171,171,170,171,171,171,171,170,171,171,171,171,171,171,171,172,171,171,171,172,172,171,171,171,171,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,171,172,172,172,172,172,172,172,172,172,172,172,172,171,171,172,172,172,172,172,172,172,172,172,172,172,174,173,173,172,170,168,171,180,192,177,187,171,178,114,188,140,175,179,154,137,180,121,160,156,169,150,122,86,176,96,176,221,182,209,139,115,133,153,191,118,48,101,175,172,162,176,164,135,77,113,135,117,112,81,167,98,142,158,182,
165,166,166,166,166,166,167,167,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,167,168,168,167,167,168,168,168,168,168,168,168,168,167,168,168,168,168,168,168,168,168,169,169,169,169,169,169,168,168,169,168,168,168,169,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,171,172,171,172,171,171,172,172,171,172,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,172,172,172,172,172,172,173,173,172,172,173,173,173,173,173,172,172,172,172,172,172,172,173,172,172,172,172,172,172,172,172,173,173,172,172,172,172,172,172,172,172,171,168,158,178,186,183,165,156,143,169,131,125,139,175,173,109,113,147,114,153,161,88,165,194,159,141,190,145,130,130,120,123,87,144,144,162,139,161,155,149,163,193,146,157,186,185,156,98,109,154,161,122,152,142,89,
166,166,166,166,167,167,167,167,167,168,167,167,168,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,168,168,169,169,168,168,169,168,169,169,169,169,169,169,169,169,170,169,169,169,169,169,169,170,169,169,169,169,169,169,169,169,169,170,170,169,169,170,169,169,170,170,170,170,170,171,171,171,171,171,171,171,172,171,172,171,171,171,171,171,171,172,172,172,172,171,172,172,172,172,172,172,172,172,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,172,172,172,172,173,173,173,173,173,173,173,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,172,173,173,173,173,173,173,174,174,173,173,173,173,173,173,173,172,99,176,179,146,186,137,166,183,126,144,158,157,134,125,156,146,155,175,110,170,130,143,187,241,184,190,149,131,137,128,169,177,157,152,188,60,106,189,204,176,167,156,131,117,151,179,163,130,175,183,131,142,130,
167,167,167,167,167,168,167,168,168,167,168,168,168,168,168,168,168,168,168,169,169,169,169,169,168,168,169,169,168,168,168,169,169,168,168,168,169,168,168,169,169,169,168,169,168,169,169,169,169,169,169,169,169,169,168,169,170,169,169,169,169,169,169,169,170,170,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,172,172,173,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,172,173,174,173,174,173,174,173,173,174,173,173,174,173,173,173,173,174,174,174,173,174,174,173,156,157,176,172,177,183,155,175,175,197,162,175,122,153,159,202,177,165,153,136,141,198,99,109,106,109,135,145,151,162,170,156,153,170,182,116,167,163,111,101,187,201,99,153,113,171,177,159,175,149,139,138,152,173,98,166,140,
167,168,168,168,168,168,169,168,169,169,168,169,168,169,169,169,169,169,169,169,169,169,169,168,169,169,169,169,169,169,169,169,169,169,169,170,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,171,170,170,170,170,170,171,170,171,171,171,170,171,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,173,172,173,173,173,173,173,173,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,173,173,173,174,174,174,174,174,173,174,174,174,174,174,174,174,174,174,174,174,175,174,174,174,174,174,175,174,174,174,174,174,174,174,174,174,174,173,174,174,174,174,175,175,175,174,174,175,175,175,175,175,174,174,175,175,175,175,175,175,177,175,176,179,162,153,172,150,182,175,183,158,207,121,158,155,205,166,178,184,141,131,191,85,149,86,119,197,148,149,147,165,115,121,139,152,119,143,144,153,127,193,174,177,165,176,161,129,146,121,197,203,135,101,137,159,94,185,
168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,170,170,170,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,169,170,169,169,170,170,170,170,170,170,170,170,171,170,170,170,170,170,170,170,170,171,170,170,170,171,171,171,170,171,171,171,171,171,171,171,171,171,171,171,171,171,170,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,173,172,172,173,173,173,173,173,172,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,173,173,173,173,173,173,174,174,174,174,173,174,174,174,174,174,174,174,174,174,175,174,174,175,174,174,174,174,175,174,174,175,174,175,175,175,175,175,174,174,173,175,175,174,175,175,175,174,175,174,174,175,175,175,175,175,175,175,175,175,175,175,176,176,175,176,176,175,175,175,175,176,176,176,178,181,167,173,171,172,170,125,141,163,131,158,134,120,149,142,149,176,118,166,117,149,175,110,138,124,94,157,107,181,116,175,196,146,113,128,194,156,182,151,168,173,190,191,166,177,142,183,112,103,118,146,140,177,169,185,187,178,126,140,
168,169,169,169,169,169,168,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,170,171,170,170,170,170,170,170,170,170,170,171,171,171,171,171,170,171,170,170,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,171,171,171,172,172,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,173,173,174,173,173,173,173,174,174,174,174,173,173,174,174,174,174,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,174,175,175,175,175,174,174,175,175,175,175,175,175,175,175,175,175,175,174,175,175,175,175,175,175,175,175,175,176,175,175,175,175,175,175,175,176,175,175,175,176,176,176,175,176,175,175,176,176,176,176,176,176,176,176,175,175,176,176,176,176,176,178,176,181,157,136,177,143,166,200,165,155,124,160,173,94,159,190,192,176,122,144,140,127,95,134,158,44,157,212,151,118,176,113,170,154,145,182,157,192,166,75,197,83,98,184,147,139,186,143,160,153,191,153,157,120,103,205,192,108,110,
169,170,169,169,170,170,169,169,170,170,170,170,170,170,170,170,170,170,171,171,170,170,171,170,170,171,171,171,171,171,171,171,171,171,171,170,171,171,171,171,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,174,174,173,174,174,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,175,175,175,176,175,176,176,174,175,176,176,175,175,176,176,176,176,176,175,176,176,176,176,176,176,176,176,176,176,177,177,177,177,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,179,178,173,216,138,156,80,148,145,171,113,150,125,159,152,88,170,149,88,186,162,161,192,152,93,157,132,93,204,159,211,187,178,154,173,147,124,163,89,90,185,148,196,186,169,138,127,161,154,102,92,174,170,185,148,125,202,161,
170,170,170,170,170,170,170,170,170,170,170,171,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,171,171,172,172,172,171,172,172,172,173,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,172,173,173,173,173,173,173,173,173,173,173,173,173,174,173,173,174,174,174,173,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,175,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,177,176,177,177,177,176,177,177,177,177,176,177,176,177,177,177,177,177,177,177,177,176,178,177,177,177,178,178,178,177,178,178,177,178,178,178,177,178,178,180,184,184,174,168,162,168,118,180,141,167,161,146,128,181,129,155,144,153,169,112,57,165,80,120,201,170,139,132,129,225,221,189,194,182,62,179,127,144,106,185,92,173,141,118,140,184,130,130,172,175,126,141,189,170,132,134,119,
170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,172,171,171,171,171,171,171,171,171,171,172,172,171,172,172,172,171,171,171,172,171,172,172,172,171,172,171,172,171,172,172,171,171,172,172,172,172,172,172,172,172,172,172,173,172,172,172,173,173,173,173,174,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,173,175,174,174,174,174,175,175,175,175,175,175,175,176,176,175,175,175,175,175,175,175,176,176,176,175,176,176,175,176,176,175,176,176,176,176,176,175,175,176,176,176,176,176,175,176,176,177,176,176,177,176,176,176,177,177,177,177,177,177,176,177,177,177,177,177,178,178,177,177,177,177,177,177,177,177,177,177,177,177,178,178,177,178,178,178,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,176,179,143,170,132,170,143,148,127,163,164,119,133,135,123,158,162,91,154,170,177,161,174,136,120,133,138,148,126,197,153,199,130,87,147,156,167,169,235,148,145,133,189,144,161,161,136,121,149,130,162,158,118,104,150,106,
170,171,171,171,171,171,172,172,172,171,172,171,172,172,172,172,171,172,172,172,172,172,172,172,172,172,172,173,173,172,172,172,172,172,172,173,172,172,172,172,173,172,172,173,173,172,172,172,172,173,172,173,173,173,173,173,173,173,173,174,173,173,173,173,173,173,173,174,173,174,173,173,174,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,174,175,174,176,175,175,176,175,176,176,175,175,176,176,177,176,176,175,176,176,176,176,177,176,176,177,177,177,176,177,177,177,177,176,177,177,177,177,176,177,177,177,177,177,177,177,177,178,177,177,177,177,178,178,177,177,178,178,177,176,177,177,177,178,177,178,178,178,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,180,178,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,178,112,173,146,155,179,117,151,177,163,107,106,155,169,153,174,132,180,113,118,180,220,170,185,140,146,160,135,172,186,152,134,183,61,89,170,154,138,199,161,161,94,125,169,157,125,100,154,145,173,157,174,167,136,176,208,
171,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,173,174,173,174,173,173,174,174,174,174,174,175,174,174,175,175,175,175,174,174,175,175,175,175,174,174,174,175,175,175,175,175,175,175,176,176,176,176,176,175,176,176,177,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,178,177,177,177,177,177,177,178,178,178,178,178,177,178,178,178,177,178,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,178,179,179,178,179,179,179,178,178,178,178,179,179,179,178,179,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,180,179,180,180,178,165,183,137,179,119,161,176,149,162,144,150,135,182,158,140,153,153,164,189,116,120,115,114,145,129,146,149,152,125,162,159,154,109,163,168,119,71,178,167,77,136,93,175,170,61,109,134,141,157,139,119,155,218,183,163,129,138,120,148,
172,172,172,173,172,173,172,173,173,173,173,173,173,173,173,173,175,173,173,173,173,173,174,174,173,174,173,174,174,174,174,174,173,173,173,174,174,173,174,174,174,173,173,174,174,173,174,174,174,173,174,173,173,174,174,174,174,174,175,174,173,174,174,175,174,175,175,176,175,174,176,175,176,176,176,175,175,176,176,176,175,175,175,175,175,176,175,176,175,175,176,176,176,177,176,177,177,177,178,177,177,177,177,177,177,177,177,177,178,177,178,178,178,177,178,178,178,178,178,178,178,178,178,178,177,178,178,178,178,178,179,179,179,179,178,177,178,178,178,179,178,179,179,179,179,179,178,179,179,178,179,178,179,179,179,179,179,179,179,179,179,179,179,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,180,180,179,180,180,180,180,180,180,180,179,180,180,180,180,180,180,179,224,109,196,92,136,179,177,170,126,194,136,183,159,105,165,170,166,177,77,163,69,116,169,120,144,118,156,111,143,149,151,110,130,148,129,143,178,130,158,142,172,160,93,132,110,175,134,149,120,147,146,131,181,160,113,156,140,119,
173,173,173,173,173,173,173,173,174,174,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,178,179,179,179,179,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,179,179,179,179,180,179,180,180,180,180,179,179,180,179,180,180,180,180,180,180,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,184,182,194,166,169,174,187,175,159,149,162,195,178,161,163,126,133,112,171,89,114,90,153,81,157,107,140,165,139,104,129,187,141,150,171,160,144,191,173,155,166,121,163,100,92,124,122,120,141,144,145,152,96,191,168,178,161,104,182,144,
173,173,173,174,173,174,174,174,174,175,174,174,175,174,175,174,174,174,174,174,174,174,175,174,174,174,175,174,175,175,175,175,175,175,175,175,175,175,175,176,176,175,175,175,174,175,175,175,175,175,176,176,175,175,176,175,176,176,176,176,176,175,177,176,176,176,176,176,176,176,177,176,176,176,177,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,179,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,179,179,179,179,180,180,180,179,179,179,179,180,180,180,180,179,180,180,179,180,180,180,180,180,180,180,180,180,180,180,181,180,180,181,180,181,180,180,180,180,180,180,180,180,180,181,180,180,181,180,181,180,180,180,180,181,180,181,181,181,181,181,181,181,181,181,182,182,182,181,178,146,159,175,152,108,223,175,98,142,146,150,124,168,147,85,130,158,139,174,80,167,199,137,92,146,100,128,130,144,163,124,168,153,59,159,78,71,169,146,127,164,137,151,115,176,120,129,119,119,187,181,179,145,85,119,156,122,183,
174,174,174,174,174,174,174,174,175,175,175,176,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,175,175,175,176,176,176,175,176,176,175,176,176,176,176,176,175,175,175,175,176,175,176,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,176,176,177,176,176,177,177,177,177,177,177,177,177,177,177,177,178,177,177,177,178,177,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,179,180,180,180,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,180,180,180,180,180,180,180,180,180,180,180,179,181,180,180,180,180,180,180,180,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,181,182,179,182,182,182,183,182,181,187,177,191,161,169,150,176,176,93,179,132,171,169,147,166,144,145,169,160,52,149,135,114,184,117,172,153,156,147,146,120,107,126,89,98,169,143,178,169,152,145,142,126,137,89,82,136,125,187,147,122,167,170,149,121,144,153,157,
174,175,175,175,174,175,175,175,175,175,174,175,176,176,175,176,176,176,175,175,176,176,176,175,176,176,176,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,176,176,176,177,176,177,177,177,177,177,177,177,177,177,178,178,177,178,178,178,177,178,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,179,179,179,180,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,180,181,181,181,181,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,181,182,182,182,182,182,182,183,182,182,182,182,182,182,173,183,169,130,174,160,149,149,217,183,180,172,189,129,138,160,173,169,156,122,97,182,166,128,100,119,107,181,106,148,104,171,183,133,169,143,54,161,117,113,93,186,67,174,128,112,137,151,122,115,166,161,123,127,167,150,119,130,95,109,189,161,130,106,
175,175,175,175,175,176,176,176,176,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,177,176,176,177,177,176,176,177,177,176,176,177,177,177,177,177,177,177,177,177,178,178,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,178,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,181,182,182,182,182,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,182,182,183,183,183,183,183,182,178,182,180,176,127,187,117,134,148,200,178,188,186,186,188,172,141,135,147,170,206,157,152,192,121,131,148,166,138,157,147,162,159,154,110,109,139,139,146,156,226,137,100,111,187,142,162,147,112,108,119,106,155,107,106,98,150,103,176,203,133,138,146,
176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,176,177,176,177,177,177,176,177,176,176,177,176,176,177,177,177,177,178,178,177,177,177,178,177,177,177,177,177,178,177,177,177,177,178,178,178,178,178,178,178,177,177,177,178,178,178,178,178,179,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,179,179,180,180,180,180,180,180,180,180,180,180,181,180,180,181,180,181,181,180,181,181,181,180,181,181,181,181,181,181,181,181,181,181,182,181,181,182,181,181,181,182,181,182,182,182,182,182,181,181,182,182,182,182,182,182,182,182,182,181,183,182,181,182,182,182,182,183,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,182,183,182,183,182,183,183,183,183,183,184,183,183,183,184,182,184,184,185,183,187,182,183,139,145,157,90,165,178,168,180,194,164,162,183,168,140,153,176,92,161,172,105,98,75,126,99,129,173,147,97,53,129,115,87,98,72,67,74,159,125,231,104,142,95,134,150,136,132,73,144,135,158,137,199,161,126,159,192,135,194,117,70,172,
176,176,176,176,176,176,176,177,176,176,177,177,176,176,177,176,177,177,177,177,177,178,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,179,179,179,180,180,180,180,180,181,180,180,180,180,180,181,180,180,181,181,181,181,181,181,181,181,181,181,181,181,182,181,181,181,181,181,181,182,182,182,182,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,182,182,182,182,182,182,183,182,183,183,182,182,183,183,183,183,183,183,183,183,183,183,182,183,183,182,183,183,183,183,183,183,183,184,183,183,183,184,183,183,184,184,183,183,184,184,183,183,184,186,184,184,47,183,183,183,185,194,83,190,166,184,158,135,135,110,133,159,99,154,150,148,161,188,90,93,96,117,110,127,187,138,129,177,132,78,164,81,126,84,134,172,181,58,77,228,108,102,112,153,121,120,139,113,113,137,215,171,177,127,134,94,118,117,137,168,90,148,
176,177,177,177,177,177,178,176,177,177,177,177,178,178,178,177,177,178,177,178,178,178,178,178,178,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,179,179,179,179,178,178,178,179,179,179,179,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,179,180,179,180,180,180,180,180,180,180,180,180,180,180,180,181,180,180,181,181,181,181,181,181,181,181,180,181,182,181,181,182,182,181,181,182,182,182,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,182,183,183,183,183,182,182,183,183,183,183,183,183,183,183,183,182,183,184,183,183,183,183,183,183,183,183,183,183,184,183,184,184,184,184,184,184,184,184,183,184,184,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,188,184,182,185,188,152,181,185,138,186,187,188,186,172,133,131,177,190,169,84,188,153,166,148,150,156,180,175,136,189,167,141,113,117,142,94,112,117,137,132,173,113,87,124,104,144,95,195,165,96,131,89,170,160,181,86,93,132,120,88,140,139,145,180,169,125,152,128,96,98,114,143,75,110,
177,177,178,177,177,178,177,178,178,177,178,178,178,178,178,178,178,178,179,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,181,180,180,180,181,181,181,181,181,181,181,180,181,181,181,181,181,181,181,181,182,182,182,182,181,182,182,182,182,182,183,182,182,182,182,182,182,182,183,182,183,183,183,182,183,183,183,183,183,183,183,184,183,183,183,183,183,184,183,183,183,183,183,184,184,184,184,183,184,184,183,184,184,184,184,184,183,184,183,183,184,184,184,184,184,184,184,184,184,185,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,184,185,217,159,145,185,199,182,181,184,187,191,162,156,160,112,151,192,216,153,163,100,186,142,185,175,221,140,167,167,185,185,161,167,125,123,139,112,115,140,150,196,142,66,100,164,117,150,155,144,118,149,77,155,113,124,168,180,134,142,131,71,133,115,190,163,168,146,83,168,131,159,90,180,111,96,
178,178,178,178,178,178,178,178,178,178,179,178,178,179,178,178,178,178,179,178,178,179,179,179,179,178,178,179,178,179,178,179,179,179,179,179,179,180,180,180,179,180,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,180,181,181,181,181,181,180,182,180,181,181,181,182,181,181,181,182,181,182,181,182,182,182,182,182,182,182,182,182,182,182,183,183,182,182,182,182,182,182,183,183,183,183,183,183,183,182,183,183,183,183,183,183,183,184,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,184,184,185,184,185,184,185,184,184,185,184,184,184,185,184,184,184,184,185,184,185,185,185,185,185,186,187,220,158,140,185,172,167,186,187,184,174,180,161,185,125,147,169,163,119,130,152,148,198,178,134,134,126,171,171,114,135,143,100,188,126,154,110,132,116,141,126,178,34,121,156,140,76,161,134,141,95,142,101,68,157,122,115,161,140,134,149,99,169,161,125,106,124,114,105,175,101,117,169,130,218,
178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,181,182,182,182,181,182,182,182,182,182,183,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,184,184,185,184,185,185,185,185,185,185,185,185,185,185,185,185,185,186,185,185,185,185,185,186,186,185,185,185,186,186,186,186,185,186,186,186,186,186,245,93,128,138,186,182,175,136,189,176,180,210,184,172,149,152,139,147,159,103,155,169,179,175,173,121,202,134,177,159,107,188,115,104,197,130,94,168,109,157,103,66,98,134,118,178,77,126,93,148,88,165,115,153,125,98,131,181,128,162,145,142,233,124,146,114,104,112,129,118,140,87,126,118,84,
179,179,179,179,179,179,179,180,180,179,179,179,179,179,180,179,179,179,179,179,180,179,179,179,179,179,180,180,179,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,180,181,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,182,183,183,183,183,183,183,183,184,184,184,183,184,184,183,184,184,184,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,184,185,185,184,185,185,185,185,185,185,185,185,184,185,185,185,185,185,185,185,185,186,185,185,185,186,185,186,185,185,185,186,186,186,186,185,186,186,185,186,186,185,186,186,186,187,186,186,186,186,186,186,186,187,187,186,187,186,186,246,115,141,187,183,160,117,180,82,188,167,99,169,150,161,177,172,142,153,147,138,196,175,136,112,89,140,143,144,157,138,114,116,84,128,123,140,121,111,158,162,94,138,149,186,94,117,142,121,123,62,90,189,179,139,150,76,188,155,113,99,111,116,122,154,170,115,141,95,48,109,104,64,169,135,
179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,181,181,182,181,182,181,181,181,182,182,182,182,183,182,182,182,182,183,183,183,182,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,185,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,184,185,185,185,185,185,185,185,185,185,185,185,186,185,185,185,185,185,185,185,185,186,186,186,185,186,186,186,185,186,185,185,186,186,186,186,186,186,186,186,187,186,186,186,187,186,186,187,187,187,187,186,187,187,186,187,186,187,187,186,187,187,187,187,187,187,187,190,86,73,152,187,189,159,141,145,185,146,150,183,185,198,144,96,111,88,96,155,178,158,155,114,170,124,137,140,157,118,150,92,192,82,132,101,87,113,88,88,164,61,75,129,185,127,150,71,105,158,188,182,172,94,137,120,150,176,63,82,79,158,167,124,184,173,164,223,157,84,190,130,82,157,164,
180,180,180,180,180,181,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,180,180,180,180,180,180,180,181,181,181,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,181,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,184,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,183,184,184,184,184,185,185,185,184,184,185,184,185,184,184,185,185,185,185,185,184,185,185,185,186,185,185,185,185,185,186,186,186,186,186,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,187,186,186,186,186,186,186,187,187,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,188,187,187,188,187,187,187,188,187,187,187,188,188,188,188,191,129,155,189,191,109,189,123,198,170,167,177,141,124,161,108,117,156,149,213,138,126,134,142,194,100,184,115,155,149,126,87,213,136,81,93,125,110,196,94,72,100,185,191,70,77,94,133,129,172,121,147,190,141,140,166,83,136,143,58,129,151,120,149,141,118,146,114,158,153,199,118,68,193,135,
180,181,181,181,182,181,181,181,181,182,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,182,183,183,183,183,182,183,183,183,183,184,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,184,185,185,185,186,185,186,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,186,187,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,187,187,187,187,187,187,187,187,188,188,188,188,188,187,188,188,188,188,188,188,188,188,188,188,189,190,125,158,190,185,187,185,121,176,163,131,187,150,171,153,143,147,148,125,141,132,175,152,116,95,163,114,125,109,205,125,184,123,184,103,122,156,138,106,150,81,165,66,180,163,161,178,107,130,209,115,145,152,102,160,153,229,113,107,70,66,103,107,172,130,212,96,120,151,229,75,110,89,141,150,
181,181,181,182,182,182,181,182,182,181,182,182,182,182,182,182,182,182,182,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,183,182,182,182,182,182,183,182,183,182,183,183,183,183,183,182,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,186,184,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,186,186,186,187,187,187,187,187,187,186,186,186,186,187,187,187,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,187,188,188,188,188,188,188,188,188,188,188,188,189,188,188,188,189,188,189,189,189,189,189,189,189,189,189,189,191,189,126,161,170,182,156,175,166,172,192,145,184,172,156,179,171,157,167,144,120,172,179,147,161,82,159,139,155,102,152,158,131,121,84,128,144,187,185,139,134,98,132,127,182,202,71,162,127,129,137,146,91,119,164,181,144,83,173,172,77,42,169,93,156,157,174,91,104,215,156,143,122,49,162,175,
182,181,182,183,183,183,182,183,183,183,183,183,183,182,183,183,183,183,183,183,182,182,182,181,182,182,182,182,182,181,182,182,182,182,182,182,183,183,183,183,183,183,183,182,183,183,183,183,183,183,183,183,184,184,184,183,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,186,186,185,186,186,186,186,187,186,186,186,186,186,187,187,186,186,186,186,186,187,186,187,187,187,187,187,187,188,187,187,187,187,187,187,187,187,187,187,188,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,187,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,188,148,133,163,192,210,195,178,178,152,153,167,165,159,194,178,183,139,158,165,152,103,213,165,168,172,186,197,138,109,84,142,109,155,85,113,150,201,91,121,86,88,98,179,161,138,168,92,189,147,97,137,129,143,154,169,125,210,158,189,177,101,178,208,182,174,61,140,132,140,116,159,155,197,93,144,
182,183,183,183,183,183,183,183,183,183,184,184,183,183,183,184,184,183,183,183,182,183,183,182,183,182,182,182,182,181,182,182,183,183,183,184,184,184,184,184,184,184,185,184,184,184,184,184,184,185,184,184,184,184,185,184,184,184,184,185,184,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,186,186,186,188,187,187,187,187,187,188,187,187,187,187,187,187,187,187,187,187,187,188,187,188,188,187,188,188,187,187,188,188,188,188,188,188,188,188,188,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,190,190,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,190,192,172,143,163,190,126,138,191,164,165,167,128,169,144,142,138,153,153,165,120,132,182,113,136,124,168,106,111,157,142,74,118,138,148,153,145,174,149,149,95,132,134,154,165,86,118,74,103,150,158,137,73,134,158,139,136,100,220,184,62,109,109,95,101,104,162,184,116,117,121,145,214,127,98,157,155,
183,183,183,183,183,184,184,184,184,184,184,184,184,184,185,184,184,184,184,184,184,183,184,183,183,182,182,183,182,183,183,182,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,185,185,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,187,187,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,190,191,191,191,191,191,191,192,191,191,191,188,174,171,163,188,194,189,171,117,125,194,194,163,184,193,174,134,167,192,152,175,155,145,160,141,137,123,121,117,132,134,103,112,146,147,123,168,155,207,170,107,144,107,76,110,79,139,157,108,191,142,48,76,102,148,156,74,95,67,106,121,103,170,84,166,143,101,168,196,98,222,155,117,108,130,122,
183,183,183,181,185,180,184,185,182,184,184,185,187,185,184,184,184,187,183,186,186,181,184,184,183,183,182,181,182,183,183,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,187,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,186,187,187,187,188,187,188,187,188,188,188,188,188,188,188,188,188,189,188,188,189,189,188,189,189,188,188,188,188,189,189,189,189,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,188,189,189,189,188,188,188,188,188,188,188,188,188,188,188,189,188,188,188,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,191,190,190,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,192,191,191,192,191,192,193,176,205,156,191,110,190,133,163,159,163,141,181,161,185,148,194,100,189,100,136,138,142,140,182,119,169,147,147,168,92,153,105,112,154,154,194,65,221,96,61,93,126,198,116,98,72,158,120,165,105,107,143,114,89,72,99,194,155,171,124,161,92,64,190,92,175,185,185,78,81,77,165,113,139,126,
171,181,180,182,184,182,182,185,177,184,184,179,187,185,163,184,187,170,185,186,169,185,186,184,184,183,182,185,182,183,183,184,184,184,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,186,187,187,187,188,188,187,187,188,188,188,188,188,188,188,188,188,188,188,189,189,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,189,189,189,190,189,190,190,190,189,190,189,189,189,189,189,189,189,189,189,189,189,189,189,188,188,188,188,188,188,188,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,192,192,192,191,192,191,191,192,192,192,192,192,192,192,192,192,192,192,192,191,212,171,162,167,188,195,158,182,179,169,174,207,172,177,153,168,187,109,159,175,130,161,155,118,91,163,159,124,101,130,97,149,226,176,177,172,69,172,122,154,92,158,155,145,194,149,112,103,148,130,180,169,60,76,81,142,86,114,134,163,93,136,186,173,159,158,167,180,70,90,109,150,101,127,79,
126,50,95,102,93,83,90,99,91,80,77,75,110,81,76,147,129,74,150,136,57,154,147,31,121,180,166,60,182,182,183,183,184,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,187,186,187,186,187,187,187,187,187,187,188,187,187,187,187,187,188,188,188,188,188,188,188,188,188,189,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,189,190,189,189,190,190,190,190,190,190,191,190,190,190,190,190,190,190,190,189,190,189,189,189,189,189,189,189,189,189,189,188,188,188,189,189,189,188,189,189,189,189,189,190,189,190,190,190,190,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,193,192,192,192,192,192,193,193,193,193,194,193,194,254,194,185,196,197,155,169,150,130,193,164,189,161,187,159,164,111,137,146,159,133,162,135,109,96,158,139,101,68,110,73,92,92,77,195,92,121,118,100,125,185,114,150,117,140,176,170,141,98,139,123,154,130,89,116,115,103,159,103,122,56,125,143,164,160,92,181,75,49,96,112,138,164,118,173,
25,29,34,26,32,101,67,122,107,82,140,108,93,120,94,102,104,92,118,98,69,150,98,61,120,11,57,30,181,182,183,183,184,185,185,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,188,187,188,188,188,188,188,188,188,188,188,189,189,188,189,188,188,189,189,189,189,189,189,189,190,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,192,191,191,191,191,190,191,191,191,191,191,190,190,190,190,190,190,190,190,190,190,189,189,189,189,189,189,189,188,189,189,189,189,189,189,189,189,190,190,190,191,190,191,191,191,191,191,191,191,192,192,192,192,192,192,192,193,193,192,192,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,190,195,241,225,89,108,136,126,186,124,180,165,155,191,165,151,136,179,161,135,133,170,149,121,198,152,129,150,140,144,101,111,191,93,109,96,135,180,84,175,65,74,139,110,168,111,135,156,156,183,142,71,201,106,104,102,211,145,110,79,113,96,160,167,171,180,86,95,178,160,114,128,93,130,146,147,58,107,
34,68,45,34,91,81,70,132,95,110,113,92,104,101,96,112,110,93,129,104,78,113,87,90,37,79,65,43,179,182,183,184,184,185,186,186,186,187,186,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,189,188,189,188,189,189,189,189,190,189,189,189,189,189,189,189,190,190,189,190,191,190,190,190,190,190,190,190,190,190,190,189,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,191,192,192,192,192,191,191,191,191,191,191,190,191,191,191,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,191,191,191,191,191,192,192,192,192,192,192,192,193,193,193,193,192,193,194,193,193,193,193,194,194,194,194,194,194,194,194,194,194,194,195,196,210,235,179,104,82,84,79,190,126,173,201,159,187,174,117,164,175,150,189,147,167,185,150,168,141,168,128,156,107,124,153,113,75,78,114,130,181,120,147,164,86,71,92,195,45,155,133,191,125,161,182,108,191,134,139,118,137,142,106,134,69,214,79,131,97,142,118,99,168,132,77,122,107,39,108,113,88,
96,75,69,130,80,45,143,80,52,149,95,64,146,112,59,139,121,67,109,146,103,74,66,139,53,69,27,50,137,182,183,184,185,185,186,186,187,187,187,188,188,188,188,188,188,188,188,189,189,189,189,188,189,189,189,189,189,189,189,189,189,189,189,190,190,189,190,190,190,190,191,191,190,191,190,190,191,190,191,191,191,191,191,191,191,191,191,191,192,190,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,193,192,192,192,192,192,192,191,191,192,191,191,191,191,191,191,191,191,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,191,191,191,192,192,191,192,192,192,192,193,193,193,193,193,193,193,193,194,194,194,195,195,195,195,195,195,195,195,195,194,195,195,195,195,195,191,239,192,252,176,142,93,94,154,164,183,196,197,168,190,167,105,174,174,182,118,153,116,170,157,127,127,183,122,80,133,179,145,169,99,158,77,166,76,188,72,110,149,141,158,128,190,152,189,128,165,219,147,187,115,187,136,138,104,107,114,71,45,148,68,168,89,158,176,169,96,72,164,146,87,114,171,120,
95,93,94,83,75,96,83,101,114,107,62,83,111,65,83,69,83,61,76,98,104,54,175,4,48,69,13,18,38,181,183,184,185,185,186,187,187,188,188,189,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,190,190,190,190,189,190,190,190,190,190,190,190,191,191,191,190,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,191,191,191,191,191,191,191,192,192,191,191,192,192,193,193,193,193,193,193,193,193,193,193,192,192,192,192,192,192,192,192,191,192,191,191,191,190,191,190,189,189,189,189,189,189,188,188,188,189,189,189,189,190,190,191,191,191,192,192,192,192,193,193,193,194,194,193,194,195,195,195,195,195,195,196,195,195,196,195,195,196,197,196,195,195,196,195,196,196,195,231,162,248,250,163,171,175,162,142,176,182,197,165,194,193,129,119,170,114,159,213,153,164,211,129,126,142,110,167,160,176,210,193,186,62,99,105,89,156,43,80,72,132,172,249,126,64,149,124,163,211,171,49,113,117,176,129,124,104,136,146,128,90,83,157,95,47,81,98,100,122,89,155,115,50,140,162,107,
113,89,99,88,105,70,72,125,85,92,132,87,86,125,83,61,159,95,57,138,142,107,23,66,73,12,12,17,25,181,183,184,185,187,187,187,189,188,189,189,189,189,190,189,189,189,189,190,190,189,190,190,189,191,191,191,191,191,190,191,191,190,190,191,191,192,192,192,192,192,193,191,192,192,192,192,192,192,193,192,192,192,192,192,192,192,193,192,192,192,192,192,192,192,192,192,192,192,192,193,193,193,193,193,193,194,194,193,193,193,193,193,193,193,192,192,192,192,192,192,191,192,192,191,191,191,190,190,189,189,189,188,188,188,188,188,188,189,189,189,190,190,191,191,192,192,193,192,192,193,193,195,194,194,195,195,195,196,196,195,195,196,195,195,195,195,195,195,195,194,196,196,195,196,195,196,196,197,180,250,250,250,156,169,170,157,197,186,188,171,176,192,184,143,163,178,152,181,167,150,154,165,133,154,166,166,176,106,120,79,128,183,176,80,108,62,88,69,147,165,158,197,195,61,118,132,74,82,135,56,121,50,197,61,205,86,135,98,120,75,112,104,171,111,132,124,142,162,155,171,166,137,123,126,134,163,
71,133,79,59,120,105,67,123,133,60,135,118,67,133,114,73,103,77,119,86,61,87,23,63,24,13,12,12,64,184,185,184,185,186,187,188,188,189,189,189,189,190,191,190,190,191,191,191,191,190,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,193,191,193,193,193,192,193,193,193,193,193,193,192,193,193,193,193,192,174,199,186,178,192,191,192,193,193,193,193,194,193,193,194,194,194,193,194,194,194,193,193,194,194,194,194,194,194,194,194,194,193,193,193,193,192,193,192,191,191,190,190,189,189,188,188,188,188,188,188,188,188,189,189,190,190,191,191,192,193,193,193,193,194,194,195,195,195,195,195,195,195,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,195,196,196,197,252,202,250,252,250,176,178,174,171,172,176,113,156,181,136,174,164,119,147,173,174,174,149,139,106,173,126,129,167,179,155,182,225,127,195,234,110,81,69,65,127,71,172,192,195,90,78,192,143,178,141,91,146,38,87,73,162,153,170,139,120,144,124,88,144,130,142,109,135,207,138,67,103,121,147,131,221,135,122,
110,73,48,110,100,66,84,115,60,67,88,123,84,65,54,111,68,56,64,94,98,13,54,75,13,12,13,11,40,89,183,184,186,187,187,189,189,189,189,190,191,191,190,190,191,191,191,192,191,191,192,191,192,191,192,192,192,192,192,192,193,193,193,193,193,193,193,193,189,194,194,193,193,194,194,194,193,193,193,194,193,194,194,194,193,106,110,105,116,84,193,193,193,193,194,193,194,194,194,194,194,194,194,195,195,194,195,194,195,195,194,194,195,194,194,194,194,194,194,194,194,192,193,192,191,191,191,190,189,188,188,187,187,186,186,187,188,188,189,189,190,190,191,191,192,193,193,194,194,194,195,195,195,195,195,196,196,196,196,196,196,196,196,197,197,197,197,196,196,196,197,197,197,196,197,197,215,247,206,242,252,250,154,175,169,165,171,180,126,181,187,149,167,121,185,112,181,121,172,173,169,115,107,164,157,167,146,135,92,110,129,141,119,82,145,162,90,166,67,75,174,162,209,117,168,92,89,78,105,158,121,74,60,96,74,122,143,150,70,104,137,93,93,136,113,70,153,118,76,80,50,117,136,88,213,124,
88,100,85,127,90,59,102,108,75,140,113,90,109,55,123,122,85,114,69,137,90,78,73,9,12,13,13,12,13,36,181,184,185,187,189,189,190,190,191,191,191,191,191,191,191,192,192,191,192,192,192,192,192,193,193,192,193,193,193,193,193,193,193,193,193,193,194,194,192,194,193,194,194,194,194,194,194,194,194,194,194,194,194,194,194,171,124,89,87,77,192,192,193,194,193,194,194,195,195,194,194,194,194,195,195,195,195,194,195,195,195,195,195,194,194,194,194,194,194,194,194,193,194,193,193,192,191,190,189,188,188,187,186,186,25,188,187,188,188,189,190,191,192,192,193,194,194,194,194,195,195,196,196,196,196,196,196,197,197,197,197,197,197,197,197,197,197,197,197,197,197,197,197,197,197,199,254,253,208,197,248,250,171,172,165,169,196,141,106,128,151,196,121,191,164,177,69,196,190,155,156,188,186,202,155,151,144,162,187,105,51,202,136,110,149,167,124,141,57,81,135,163,140,60,96,143,70,77,165,66,149,64,146,147,107,117,171,120,193,74,152,100,205,100,176,149,127,114,55,127,56,56,95,53,168,111,
130,94,64,116,100,97,101,87,128,82,58,138,101,76,89,104,135,102,66,51,20,65,120,16,13,14,13,13,14,51,188,184,185,188,189,190,190,190,191,191,191,191,192,192,192,192,193,192,192,193,193,193,193,193,193,193,193,193,193,193,194,194,194,194,194,193,194,194,194,192,195,194,194,195,194,194,194,194,195,194,194,194,194,194,196,175,171,175,177,102,194,192,193,194,193,194,194,195,195,194,195,195,196,196,195,196,195,195,196,195,195,195,195,195,195,195,195,195,195,194,194,194,193,194,194,192,191,190,189,188,188,186,187,25,18,48,190,189,188,189,190,191,192,192,193,194,194,195,195,195,196,196,196,196,197,197,197,197,197,198,197,197,198,197,198,198,198,198,198,198,198,197,200,199,199,201,254,238,215,126,249,250,159,170,169,166,169,129,163,120,100,185,178,123,160,157,166,187,108,169,124,162,139,122,186,112,192,157,83,155,165,99,126,151,83,119,84,111,107,69,77,198,218,56,166,143,149,157,152,105,81,141,110,221,73,106,151,70,103,34,174,176,122,89,140,166,129,121,87,62,129,112,62,69,120,101,
139,142,94,80,110,122,84,56,122,147,84,89,133,122,80,71,118,172,108,20,50,71,137,26,11,13,14,13,11,74,185,183,186,188,190,190,191,191,191,192,192,192,192,192,192,192,193,192,192,193,193,193,193,193,193,193,193,193,194,194,193,194,194,194,194,194,194,194,198,192,194,194,194,197,194,194,195,194,195,194,194,194,195,195,195,179,181,173,173,94,190,192,192,193,193,194,195,195,195,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,195,195,195,195,194,194,194,194,193,193,192,191,189,188,187,187,23,17,29,39,46,192,189,189,190,192,192,193,194,194,195,195,195,196,196,197,197,197,197,197,198,198,198,198,198,199,198,199,199,199,199,199,199,199,199,199,224,198,199,214,254,147,193,120,249,250,167,178,172,172,207,200,180,155,185,135,192,157,148,198,189,191,158,201,185,179,184,151,139,144,211,161,134,153,119,159,125,80,114,121,133,172,180,80,70,82,219,122,94,59,68,98,84,100,63,131,134,134,99,163,165,153,78,115,94,188,140,102,166,87,89,124,87,112,155,140,96,160,189,115,
121,63,80,118,75,88,59,147,112,46,110,114,103,79,42,156,111,86,39,70,68,57,145,124,8,10,9,11,10,12,38,182,186,188,190,190,191,192,191,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,194,194,194,194,194,193,184,194,194,194,194,195,195,195,195,186,195,195,195,190,195,195,196,195,197,193,195,193,197,195,194,176,182,174,173,77,190,189,189,192,190,193,195,194,196,199,198,196,195,196,196,196,197,197,197,196,198,197,197,193,197,197,195,197,198,196,193,196,192,195,191,193,191,192,189,189,188,26,22,27,26,47,35,41,190,189,193,191,193,193,193,195,195,196,196,196,197,197,197,197,198,198,199,199,199,199,199,199,199,200,200,200,200,200,200,200,200,200,205,178,200,248,255,150,197,117,250,250,152,168,170,163,205,154,170,193,179,187,121,167,171,180,143,171,106,150,185,179,161,178,136,148,154,190,119,190,201,70,114,90,156,130,165,135,202,119,54,76,55,81,113,83,97,203,85,99,176,128,127,99,229,144,113,168,99,148,165,85,125,124,169,187,216,105,95,51,120,171,59,125,176,96,
54,140,122,69,112,111,115,94,78,147,125,81,111,72,146,110,77,67,8,51,63,88,151,134,14,12,13,12,11,17,30,185,186,189,190,190,191,191,192,192,192,192,193,193,193,193,193,193,193,194,194,194,194,194,194,195,195,195,195,195,196,195,195,196,196,196,196,196,196,194,195,195,196,195,196,196,195,195,191,74,170,167,70,168,192,183,173,177,171,29,25,34,50,40,104,101,190,192,121,197,195,176,195,196,191,198,192,198,199,197,197,198,197,195,196,193,198,196,196,198,197,194,197,195,193,196,194,191,192,191,20,18,29,22,25,11,42,38,45,192,194,195,194,194,194,195,196,196,197,197,196,198,198,198,199,199,199,200,200,200,200,200,200,200,200,200,201,200,200,201,200,201,200,203,171,253,194,141,195,130,250,250,163,169,179,171,195,131,194,195,149,149,159,157,168,184,142,162,173,89,184,124,186,144,161,166,92,177,203,221,139,146,167,124,113,134,75,115,195,114,177,61,49,82,185,55,98,168,153,82,192,131,75,112,166,171,159,165,189,134,82,150,54,106,76,191,72,62,92,73,65,124,93,130,148,178,
71,75,116,118,110,74,124,124,69,91,88,133,121,85,79,102,106,71,44,74,94,93,120,141,22,11,12,12,10,10,68,187,187,188,189,191,191,192,192,193,193,193,194,194,194,194,194,194,194,195,194,195,195,195,195,196,195,196,196,195,195,195,196,197,196,197,191,196,197,196,196,196,197,199,196,197,195,195,161,162,140,118,136,120,179,186,147,170,141,14,19,27,40,35,39,42,71,151,187,86,136,164,165,114,119,96,84,140,124,117,164,142,148,166,150,105,153,132,108,151,103,125,98,88,109,136,112,164,140,20,16,27,21,12,10,6,29,41,41,51,165,84,160,171,150,178,195,185,190,200,199,200,191,199,199,199,200,200,202,202,201,198,201,201,200,203,192,203,203,179,201,202,202,202,201,187,204,210,148,164,250,250,172,173,179,171,193,157,181,170,133,182,177,128,184,123,115,125,107,112,138,187,152,102,141,86,158,128,135,184,133,133,170,135,158,113,118,72,90,157,76,118,107,84,57,190,103,160,126,160,181,149,122,67,98,168,175,151,145,198,119,140,130,131,149,167,124,89,146,194,122,156,69,139,150,97,
116,84,76,88,82,90,83,56,105,77,93,96,68,107,78,121,78,31,70,99,99,94,91,145,115,8,10,9,11,10,16,85,187,189,190,191,192,193,193,193,193,194,194,194,195,195,195,195,195,195,195,196,196,196,196,196,196,191,195,188,198,197,197,197,196,197,195,197,198,199,197,197,198,198,197,197,190,196,56,50,134,157,118,147,32,45,52,47,96,18,71,184,81,59,78,95,64,57,100,69,76,113,142,106,85,71,129,107,88,163,120,88,175,133,88,160,121,87,169,111,83,89,92,87,94,98,83,153,23,13,26,24,16,19,15,17,9,46,39,48,59,187,180,133,155,183,90,126,178,79,143,149,83,144,137,53,149,129,48,148,140,103,161,118,142,170,122,141,176,102,195,145,80,148,131,100,153,93,114,195,250,250,164,178,177,173,136,115,145,162,139,153,175,192,166,141,169,77,85,194,124,93,116,137,172,130,161,125,143,157,161,155,130,133,73,86,106,180,124,167,139,162,210,86,75,66,153,129,131,144,190,159,168,121,112,144,62,118,195,138,118,124,90,95,93,107,125,120,122,169,114,103,110,113,175,83,
106,58,134,93,71,129,134,122,82,56,135,106,115,110,90,60,17,44,80,98,99,96,92,148,126,13,7,8,10,9,17,29,187,189,191,192,193,193,193,194,194,194,195,195,195,196,196,196,196,196,196,196,196,196,197,197,197,198,197,182,194,198,194,199,198,199,197,198,198,196,181,200,197,200,198,198,190,195,10,126,92,153,149,83,92,132,128,136,158,110,35,162,107,90,144,89,99,140,79,100,130,100,102,135,93,137,171,110,138,185,125,114,159,171,87,173,157,122,196,114,133,154,122,118,150,135,97,20,16,25,22,13,22,21,17,22,13,12,51,35,50,59,160,160,113,150,164,44,69,82,69,148,97,131,135,124,155,176,125,144,181,122,170,169,119,166,112,131,148,126,99,115,122,110,151,106,149,155,123,249,250,250,151,176,173,174,167,94,136,162,128,155,201,128,111,97,167,195,174,155,126,203,126,137,196,153,123,134,159,111,107,134,82,134,138,67,134,165,106,108,135,68,234,123,65,171,173,177,108,151,191,138,194,126,151,191,82,134,195,135,135,101,71,128,72,55,77,129,150,142,131,201,82,112,151,60,
67,63,43,70,121,71,33,100,88,93,60,49,48,50,97,61,51,67,98,99,98,97,96,120,133,26,18,15,17,15,14,68,187,189,190,192,193,193,194,194,195,195,195,195,196,196,196,196,196,197,197,197,197,197,197,197,197,198,200,191,171,198,194,198,199,186,198,196,198,197,202,198,196,200,192,197,198,193,128,78,119,97,74,127,105,68,107,79,51,110,117,83,159,126,71,153,172,112,127,170,164,108,197,201,93,70,180,106,102,187,141,78,195,144,82,201,167,93,232,195,93,232,164,77,200,223,19,15,19,20,11,15,22,19,17,23,17,17,9,66,36,54,37,189,146,74,158,118,82,88,89,149,160,109,219,176,150,193,186,133,192,182,142,207,173,132,220,169,146,204,146,145,192,166,165,211,161,190,214,249,249,250,156,177,181,179,197,63,164,120,130,180,186,93,139,107,144,186,144,163,113,100,192,126,157,197,124,133,161,148,184,95,146,129,164,60,66,124,181,159,68,167,192,154,136,79,127,102,116,123,206,169,197,150,132,178,116,106,171,175,179,100,83,132,98,172,112,165,122,137,49,193,63,176,91,90,
64,131,115,123,90,35,140,120,105,95,73,70,39,140,49,22,73,95,96,99,99,99,96,89,142,35,21,21,17,17,20,28,150,190,191,192,193,194,194,194,195,196,196,196,197,197,197,197,197,197,197,197,197,199,198,198,195,197,197,200,190,199,191,199,199,200,196,194,197,196,200,198,194,200,181,198,196,96,164,113,96,142,171,87,117,180,94,71,180,174,88,202,202,107,134,192,133,93,130,180,102,150,209,139,62,198,157,84,183,188,105,121,192,133,75,192,167,116,180,168,141,131,174,98,61,21,15,23,19,11,15,18,23,21,23,25,19,17,18,4,63,37,53,42,77,82,159,172,125,188,190,137,198,190,160,203,174,201,209,190,191,212,179,150,204,185,135,214,196,156,217,188,160,206,182,166,217,205,194,249,249,247,145,175,173,168,202,70,73,193,160,136,197,123,172,137,156,140,110,110,208,162,126,167,126,230,166,109,140,223,64,114,129,97,113,93,84,106,208,45,111,107,194,95,100,101,110,140,156,173,172,193,190,107,145,101,135,68,123,88,84,60,73,121,157,76,49,42,70,61,35,45,55,85,67,95,
152,113,70,100,102,152,87,62,99,55,155,125,131,102,77,39,75,97,99,101,100,99,97,93,143,40,22,23,23,21,17,50,36,190,191,193,193,194,195,195,196,196,197,196,197,197,197,198,198,198,198,198,196,200,199,199,198,194,188,197,203,197,196,200,200,198,196,195,192,201,201,199,190,200,192,196,189,12,84,99,126,179,102,98,185,116,48,203,169,115,188,205,109,108,194,145,80,105,175,97,79,168,155,82,139,158,92,97,140,108,82,119,115,58,101,116,61,101,99,81,80,152,122,63,21,14,20,22,14,16,16,17,24,23,23,23,22,16,20,11,9,66,36,66,63,168,119,202,167,174,213,164,110,180,143,93,154,161,81,169,136,70,177,158,82,171,183,98,136,197,117,145,209,137,146,215,170,186,197,250,251,245,161,172,195,190,73,182,84,193,141,181,203,149,159,169,122,198,162,196,177,106,92,109,173,102,200,199,173,125,62,223,150,222,68,83,175,83,96,145,89,99,132,82,199,81,49,144,83,91,199,204,167,218,173,136,147,102,130,82,157,143,127,119,207,67,54,61,138,187,101,62,117,66,46,79,
97,102,94,69,72,149,146,73,78,85,77,113,97,99,65,74,98,97,98,100,99,100,97,94,119,37,18,17,20,15,36,13,49,193,191,193,194,195,195,196,196,197,197,197,197,197,198,198,198,199,199,199,199,190,199,201,201,186,187,194,196,199,203,201,201,201,201,186,201,202,203,195,188,201,200,199,187,106,80,98,179,115,68,178,140,79,152,182,115,85,156,123,66,112,122,81,76,142,109,98,104,110,55,149,103,95,81,155,118,85,187,160,114,179,194,142,160,186,156,121,150,129,99,80,16,20,19,26,17,20,20,18,23,23,22,19,21,19,16,17,20,35,58,45,56,82,132,145,177,120,88,125,87,113,151,117,128,165,137,118,183,132,75,182,144,87,170,143,110,180,167,110,112,168,124,135,148,144,204,249,249,246,174,180,178,170,15,18,17,85,183,165,175,206,183,176,132,174,209,106,160,109,43,108,150,125,110,185,132,130,113,77,105,162,98,140,198,175,57,82,129,132,107,148,97,30,82,127,106,101,164,179,172,162,96,136,205,118,145,167,219,129,75,159,175,113,116,123,99,101,109,87,93,69,63,154,
108,128,105,66,126,102,125,93,78,72,54,82,26,21,52,84,100,98,99,101,101,100,101,95,89,130,97,14,16,19,13,12,46,187,190,193,194,195,196,196,196,197,197,198,198,198,199,199,199,199,199,199,200,202,178,200,200,200,199,193,200,201,201,202,202,201,185,157,202,201,201,202,201,204,198,200,121,79,163,108,78,140,129,109,99,139,126,104,99,107,98,57,128,120,55,118,159,133,83,113,172,136,149,187,202,135,183,206,147,122,193,169,97,143,183,118,97,201,172,114,209,189,101,102,25,17,5,9,20,21,21,19,19,22,23,23,21,21,22,22,20,11,1,60,43,55,130,118,142,146,98,172,188,108,167,194,142,184,207,167,162,213,158,152,212,204,163,212,215,180,198,220,179,160,109,194,176,128,190,248,249,248,178,177,170,171,23,25,32,6,205,156,158,217,179,175,164,156,90,133,104,112,183,177,191,122,127,89,110,97,100,141,194,78,114,190,138,162,101,69,180,195,183,118,67,50,137,125,110,159,106,174,143,101,180,163,194,115,121,153,195,90,54,163,182,106,183,138,163,169,117,214,149,160,133,114,
66,99,100,113,102,69,74,61,107,164,124,61,62,33,55,79,97,100,97,100,101,100,101,97,93,143,120,9,13,12,13,11,21,44,193,193,195,195,196,196,197,198,198,198,199,199,199,200,200,200,200,201,201,201,200,200,181,203,201,194,172,199,198,196,200,204,201,177,197,186,203,204,203,198,193,200,21,200,140,75,188,160,100,164,180,119,103,124,160,95,68,184,146,85,149,169,170,79,65,198,152,79,121,184,146,87,129,175,106,66,204,160,75,186,193,98,142,202,179,102,138,193,122,116,81,6,3,14,18,21,23,20,20,19,20,22,23,22,21,19,19,6,4,7,54,44,168,140,169,206,173,158,210,155,125,200,188,100,188,191,113,140,186,145,114,208,203,129,189,216,184,166,217,170,155,184,229,231,200,252,249,248,178,173,172,178,33,31,34,15,158,159,191,142,157,172,161,168,70,194,88,91,145,126,122,147,99,159,122,115,145,135,115,106,112,72,183,192,77,62,142,141,123,145,192,112,139,153,182,110,78,163,194,171,169,170,182,201,146,114,107,70,76,107,89,70,153,174,117,181,137,168,125,177,121,115,
124,94,119,113,60,59,50,104,115,166,110,112,69,74,46,97,98,99,102,100,102,101,101,100,97,117,134,12,10,11,12,12,17,35,192,193,195,195,196,197,198,198,199,199,200,200,200,201,201,201,202,199,201,201,188,203,200,188,166,199,205,122,203,202,195,204,203,159,203,188,211,192,202,200,179,202,15,130,63,174,144,69,181,200,112,132,151,173,116,54,200,187,127,140,149,159,98,57,173,162,92,119,103,109,86,84,176,136,117,137,131,109,69,165,152,85,103,136,132,113,129,96,74,119,86,4,4,15,17,33,34,22,21,17,19,22,22,23,67,65,19,8,2,5,14,79,213,198,109,206,202,133,135,187,149,83,108,164,99,108,147,64,127,110,82,166,136,133,111,94,154,165,101,125,186,166,115,229,206,226,248,248,172,173,174,181,32,30,27,26,10,179,202,158,81,138,179,150,190,141,117,132,168,142,120,101,100,111,137,112,84,117,151,127,80,187,163,188,169,63,101,125,158,107,121,99,60,109,103,165,148,109,156,197,203,159,198,126,113,112,100,122,155,141,175,54,108,164,127,142,94,115,112,149,117,153,
91,58,92,74,148,142,103,100,80,49,21,25,37,59,98,100,98,101,101,101,102,102,102,99,96,87,139,107,8,13,13,12,12,55,193,191,194,195,197,198,199,199,199,200,200,200,201,201,201,201,202,201,203,202,205,204,205,200,151,197,208,207,207,202,198,205,197,179,197,195,141,202,201,186,191,133,98,130,135,87,75,164,158,93,72,168,153,88,69,172,150,83,57,123,129,67,83,118,99,85,129,160,89,92,165,153,110,120,153,138,114,100,182,152,74,134,171,142,108,99,169,141,108,99,93,8,2,18,18,33,32,22,22,21,25,41,25,21,66,66,21,10,3,1,9,90,55,178,99,117,68,76,88,127,117,113,88,204,148,102,199,204,170,155,192,194,146,150,206,173,149,222,184,100,181,191,154,126,157,133,245,245,166,178,180,183,27,11,23,19,9,188,138,180,161,147,166,99,186,94,131,104,184,180,121,195,139,94,88,50,149,107,70,140,154,171,141,209,196,43,133,206,125,142,94,175,64,174,122,202,184,86,132,188,198,128,158,161,158,100,78,123,133,190,133,103,44,132,199,110,118,168,172,132,121,167,
119,105,84,86,52,63,97,72,75,29,131,41,64,99,97,98,103,104,103,103,104,101,101,98,97,93,145,129,16,14,14,14,13,16,89,192,194,197,197,199,199,199,200,200,200,201,201,201,201,202,202,203,202,202,173,199,204,179,196,203,194,187,202,205,204,205,196,178,200,171,199,204,201,136,180,34,130,102,58,194,148,82,184,159,104,100,73,171,154,61,68,107,188,133,83,196,200,155,91,90,181,127,123,146,166,179,82,75,208,200,127,139,171,188,113,91,207,195,108,155,178,190,82,41,52,3,2,21,19,32,33,19,24,96,25,28,25,23,67,67,21,10,0,2,13,99,46,203,200,156,114,197,199,115,129,223,173,100,218,203,172,208,208,179,166,201,198,158,162,222,202,164,221,207,209,186,205,230,218,138,188,247,181,176,187,182,26,20,34,37,36,23,117,174,104,188,132,127,192,136,99,119,128,206,181,154,81,80,110,122,158,106,72,122,109,208,139,190,97,119,158,135,170,114,65,184,199,118,209,130,166,165,78,91,193,165,211,166,81,41,124,222,82,180,52,102,223,122,88,131,133,196,182,127,111,141,
145,114,74,78,66,76,51,122,43,49,44,56,95,99,100,100,102,99,101,104,103,102,102,98,99,94,113,134,20,14,15,14,14,23,21,193,195,197,198,198,199,200,201,201,201,201,202,201,202,202,202,202,202,203,202,205,205,206,195,188,204,150,150,191,185,199,207,198,189,170,202,206,187,191,175,24,105,84,190,139,72,193,207,125,101,71,209,163,98,121,141,184,135,60,188,198,161,86,59,185,159,74,78,151,185,137,105,117,182,175,95,81,177,185,134,103,174,184,84,84,195,190,35,73,3,4,1,72,26,21,28,20,25,24,23,26,25,21,68,68,22,12,2,1,10,17,140,52,208,203,121,172,201,203,99,111,206,175,129,162,178,147,81,146,154,94,77,150,123,93,156,179,171,91,132,227,222,182,222,216,141,242,150,169,171,79,24,31,35,35,35,3,187,169,166,188,116,165,172,149,182,156,148,132,162,128,128,131,137,100,142,85,207,142,117,185,180,106,79,106,167,166,90,183,113,160,189,165,146,132,167,186,101,104,99,205,210,99,58,109,147,139,111,171,98,91,136,70,142,61,112,182,119,167,119,79,
83,57,102,146,125,103,89,82,57,8,36,64,97,100,100,100,98,99,124,107,104,106,105,99,98,96,88,141,116,11,15,13,12,13,63,192,195,197,198,199,200,200,201,201,201,202,202,202,203,203,203,203,196,203,203,191,203,199,205,176,204,205,165,205,197,207,205,205,157,191,194,194,179,207,140,102,107,147,100,80,130,192,141,89,81,190,174,143,72,99,152,111,85,66,149,110,75,68,110,146,86,141,152,123,97,81,88,148,152,67,134,131,123,100,58,162,146,94,104,121,146,83,44,123,171,129,3,64,36,19,20,20,18,18,22,27,26,17,72,64,20,12,10,1,14,7,20,50,105,116,125,103,67,52,125,83,140,127,78,115,124,127,128,129,187,172,121,138,180,158,120,118,183,158,104,143,141,124,175,201,123,182,113,73,96,93,4,31,28,24,22,29,45,136,131,150,194,197,180,161,157,185,144,140,96,158,127,161,169,121,188,214,128,156,178,131,145,164,164,166,147,141,155,167,202,148,54,72,118,185,163,201,164,94,86,192,195,74,130,132,91,72,133,107,79,96,108,80,116,54,99,105,158,95,88,134,
64,137,95,142,116,144,136,115,56,54,61,97,96,99,99,99,157,128,99,103,103,102,101,103,99,96,92,146,128,15,16,13,13,13,20,171,196,197,198,199,200,200,201,201,202,203,203,203,203,204,204,195,207,190,201,188,205,188,202,202,189,202,204,202,205,208,206,206,154,210,193,208,189,124,38,183,114,63,187,163,97,111,97,163,155,103,90,88,180,153,119,111,112,168,147,89,154,158,177,144,164,198,167,150,103,61,202,206,147,97,89,208,192,139,126,153,194,116,74,203,216,190,85,90,221,227,11,78,36,20,22,16,20,21,23,22,18,21,19,21,20,11,1,7,13,23,23,26,27,109,188,169,143,85,206,201,175,165,204,185,147,119,214,200,163,198,215,195,151,152,208,200,141,209,226,208,187,171,227,228,147,207,199,86,163,99,56,113,125,146,114,170,71,194,135,153,211,195,186,134,124,120,133,169,228,139,100,169,129,155,195,150,155,159,156,63,151,119,157,145,149,169,203,130,183,149,144,81,81,199,136,214,216,211,128,134,178,195,165,176,125,48,86,82,139,115,97,50,131,144,57,157,86,97,61,145,
79,105,85,68,72,50,94,27,39,48,87,96,97,101,101,98,161,156,103,113,103,101,103,103,102,99,92,110,136,21,11,11,8,10,18,27,196,197,198,200,200,201,202,202,203,203,203,204,204,201,204,204,205,205,161,197,196,201,194,207,182,194,193,167,192,205,209,208,165,137,205,205,198,144,9,160,66,184,203,118,121,95,186,194,135,87,73,201,193,125,86,91,197,199,134,95,67,186,199,147,114,157,139,140,115,125,153,192,137,88,158,204,179,104,59,181,195,140,69,129,188,168,104,108,145,195,35,72,38,21,22,19,22,18,24,48,22,23,36,74,19,11,2,21,22,38,41,35,39,41,51,138,204,146,122,201,200,175,106,164,181,137,100,126,169,158,87,120,191,136,113,153,171,178,107,106,216,221,194,169,194,120,70,88,94,101,97,133,150,210,212,177,24,123,173,108,194,210,219,142,137,209,197,173,142,169,125,164,173,150,180,160,193,157,137,74,103,155,124,136,120,101,180,170,159,98,116,139,125,158,165,180,187,196,145,113,106,198,117,184,170,133,113,93,67,75,97,110,75,56,71,161,60,145,88,174,
93,45,70,80,63,21,145,135,32,61,96,93,97,100,100,100,158,103,149,162,104,128,113,98,102,100,94,90,142,121,10,8,9,9,9,51,198,197,198,200,201,202,203,202,203,204,204,204,205,204,200,207,182,199,140,190,194,199,204,208,203,212,203,181,202,187,207,210,184,192,169,198,203,124,91,104,142,173,140,71,82,183,162,105,65,42,193,174,128,94,65,123,147,116,112,100,106,93,75,57,113,84,92,83,64,104,109,80,106,84,119,132,87,76,113,122,116,75,135,146,111,99,87,169,180,137,47,69,36,20,19,17,23,20,23,44,26,17,49,69,18,11,37,19,11,26,33,23,28,32,25,16,25,148,107,103,94,102,103,52,150,149,110,117,131,216,185,115,187,200,149,134,110,212,155,102,119,140,112,137,137,127,127,136,128,85,119,128,224,181,72,164,100,98,80,121,164,217,126,165,126,205,161,214,181,121,148,167,182,134,162,183,189,98,84,180,169,130,151,107,178,82,182,139,179,141,155,152,118,72,117,183,122,186,207,157,164,179,154,214,119,116,156,92,79,148,59,88,139,62,88,123,62,83,120,122,
39,80,37,98,89,45,119,60,54,96,94,96,98,101,98,102,156,61,80,139,103,161,157,145,99,98,95,93,147,129,15,18,20,20,17,42,197,197,199,200,202,203,203,204,204,204,205,205,206,206,206,206,204,203,192,207,189,200,205,158,209,207,205,207,209,210,208,196,207,197,199,157,201,34,200,196,121,119,129,160,126,65,112,121,173,135,100,75,68,217,212,164,93,48,206,206,181,117,95,168,144,85,68,129,189,195,165,100,72,181,214,172,119,61,215,217,170,113,55,209,212,192,96,106,226,226,43,68,34,28,20,16,23,21,24,46,28,16,60,70,18,11,5,24,12,13,16,19,34,27,29,28,40,38,106,161,157,185,199,162,107,201,202,171,135,162,202,186,137,196,202,201,165,110,222,212,205,192,137,222,225,206,148,93,188,191,120,131,87,161,189,113,154,85,153,217,208,196,105,129,118,114,169,111,227,147,204,182,111,71,134,165,168,132,147,142,142,124,156,193,75,80,148,163,99,191,201,142,129,152,193,178,143,178,187,157,89,131,137,149,156,117,91,53,89,174,119,69,142,171,99,96,145,153,149,154,
83,44,118,36,40,22,14,36,46,97,95,98,100,101,100,100,158,24,85,152,101,132,135,159,109,98,96,92,112,132,22,21,21,19,19,31,51,198,200,201,203,204,204,204,204,205,206,206,207,208,209,198,206,208,150,150,204,209,207,208,207,164,180,203,140,211,208,176,150,198,204,202,174,10,194,114,125,111,183,147,114,105,122,198,191,106,77,67,195,201,159,111,80,153,176,182,129,112,108,132,159,67,96,147,122,181,173,83,101,148,198,176,143,84,92,205,179,146,65,115,198,196,119,83,91,192,51,72,32,28,30,16,20,19,52,41,27,16,73,72,16,12,60,45,18,15,28,36,31,24,35,40,39,37,43,48,73,178,198,194,119,73,204,198,176,74,66,182,168,167,71,127,208,191,155,147,177,224,211,171,196,214,224,206,192,176,158,219,202,196,162,187,193,78,97,193,165,161,160,148,95,177,175,165,108,113,125,217,109,69,124,189,179,75,112,129,116,199,165,145,108,98,141,145,90,212,171,135,184,188,82,204,167,214,210,158,108,146,76,170,196,75,145,89,52,147,55,73,124,69,69,41,97,101,145,81,
145,148,172,127,54,2,28,54,90,96,95,98,99,99,98,101,156,26,87,158,101,108,80,89,106,100,96,93,87,141,23,24,23,24,23,17,38,199,200,202,203,204,204,205,205,206,207,207,207,208,193,194,200,203,206,207,173,182,210,210,178,206,192,211,206,188,199,200,202,161,174,196,155,130,168,127,130,133,88,109,80,131,165,125,98,48,73,135,150,74,73,95,131,129,132,83,125,98,140,134,155,186,145,134,115,87,89,67,120,139,107,109,89,133,142,124,123,80,160,151,141,115,85,125,161,205,66,62,30,26,29,17,85,91,98,115,20,18,63,63,19,9,20,47,19,17,24,21,17,18,35,32,27,16,24,29,28,25,65,150,131,85,111,113,126,103,84,131,143,146,135,106,159,165,155,139,76,126,106,140,142,113,123,107,164,179,156,129,149,189,170,127,82,125,79,153,179,181,198,156,147,128,132,127,164,106,205,119,138,42,187,114,142,73,88,138,164,198,187,189,110,147,135,119,158,147,149,133,144,104,94,206,205,213,160,161,189,125,104,114,117,111,114,115,98,108,95,135,154,164,76,99,145,178,147,131,
155,124,159,63,12,56,51,59,92,99,95,99,100,100,100,101,155,23,88,159,101,94,85,94,98,97,97,96,91,143,27,23,21,20,21,8,50,197,201,203,204,205,206,206,207,207,208,207,207,208,209,207,193,197,202,205,201,147,208,207,212,197,159,208,173,209,198,175,178,216,187,205,62,156,197,114,116,56,198,194,142,106,95,143,134,193,189,146,85,56,194,174,186,111,94,105,128,198,193,139,161,187,144,186,151,110,74,169,187,188,180,109,158,173,205,180,138,97,76,216,201,173,85,107,212,222,91,76,69,87,97,91,87,95,92,74,64,39,15,15,12,7,20,31,15,14,16,15,24,28,25,29,23,34,32,41,39,35,44,43,203,207,175,140,158,207,204,181,162,147,208,203,189,158,155,213,203,198,169,130,180,196,174,156,122,154,165,184,171,141,144,158,202,181,102,80,123,159,160,114,112,77,176,198,122,97,177,155,192,120,114,191,151,156,164,179,149,135,145,177,162,186,111,197,93,153,200,162,133,146,101,178,176,115,189,133,132,192,95,122,145,89,152,152,185,203,113,94,136,57,114,51,133,172,164,132,
125,119,76,48,11,28,43,91,92,96,96,100,100,100,99,100,155,27,88,161,101,88,87,94,99,99,98,96,91,117,115,14,11,14,12,13,22,92,201,203,204,205,206,206,207,208,208,209,209,210,207,199,200,208,211,195,163,206,160,168,209,212,194,198,208,189,192,195,159,191,208,170,7,139,103,104,102,188,187,122,85,52,157,169,179,174,113,85,73,194,215,170,129,81,120,82,174,193,143,94,134,113,114,151,127,100,94,103,186,201,149,97,69,188,192,133,114,105,68,127,172,162,86,77,111,158,45,64,36,44,19,33,30,39,34,23,78,29,22,22,24,8,32,44,31,22,28,29,26,36,35,34,36,46,45,36,44,45,50,47,42,123,206,183,137,93,211,207,194,172,135,171,205,196,185,165,179,185,204,199,183,162,167,210,197,195,167,150,189,200,191,153,148,199,198,86,173,162,217,165,162,74,115,154,146,180,200,152,195,156,105,115,85,130,110,176,174,158,158,115,133,146,86,159,99,67,93,90,134,96,125,162,184,142,204,123,100,187,213,101,89,108,90,141,150,177,148,48,74,67,84,106,127,135,181,144,
135,45,132,3,31,52,93,92,94,96,100,97,101,99,102,103,155,37,87,159,100,87,88,94,101,102,97,95,93,83,131,85,10,14,14,14,18,29,203,204,205,206,207,207,208,209,209,210,210,206,206,213,206,212,206,193,205,214,203,198,181,212,204,197,209,161,205,206,214,207,214,163,90,186,178,105,109,70,117,110,165,128,123,94,71,108,86,170,159,108,101,62,145,179,136,138,103,91,56,181,107,137,75,99,129,157,168,153,121,119,72,191,171,163,138,135,99,75,217,216,191,95,61,167,193,194,167,38,52,46,16,37,36,36,55,23,97,49,24,70,34,9,18,38,31,20,23,33,19,40,11,33,29,31,46,35,19,19,33,36,36,27,48,53,143,138,114,81,99,106,91,110,103,95,85,115,127,133,147,96,136,166,164,142,88,97,188,170,142,88,83,96,92,111,115,31,110,146,202,172,206,104,132,173,218,181,145,151,239,165,44,150,154,126,190,143,199,174,77,92,108,126,218,165,174,100,51,49,148,77,77,51,94,192,84,64,129,191,127,70,75,135,81,148,88,121,167,50,31,77,44,46,124,142,141,119,
36,33,26,27,48,75,92,90,91,96,99,99,99,98,100,102,154,51,87,158,99,76,90,93,101,99,97,96,94,90,141,119,9,15,13,13,12,74,203,204,205,206,207,208,209,209,211,210,211,213,198,210,205,196,212,212,210,199,209,137,214,205,200,169,133,206,203,201,182,192,198,56,128,210,165,106,78,169,98,204,191,135,88,73,167,182,186,180,144,78,60,176,187,185,168,84,129,73,213,217,165,156,194,142,89,218,213,163,144,92,148,117,199,211,172,108,76,191,189,197,198,115,103,89,203,160,188,139,95,70,115,80,121,76,90,81,105,40,24,65,86,16,24,121,61,146,118,122,115,161,66,119,135,118,155,155,118,106,106,169,60,134,127,126,147,198,215,197,169,149,113,206,210,186,157,159,207,214,217,186,180,169,140,235,216,204,168,173,208,209,199,173,155,222,198,144,100,107,183,173,134,84,143,156,129,185,187,224,212,103,157,131,191,225,136,152,117,143,143,62,76,113,157,115,76,30,132,86,160,116,75,125,127,68,57,130,159,199,143,131,79,67,143,88,133,181,173,48,57,38,133,97,89,98,70,72,
25,20,21,53,53,90,95,93,91,96,97,99,100,101,101,100,155,49,89,159,97,68,92,95,101,100,99,97,95,89,114,128,18,12,14,11,13,21,167,204,206,207,207,209,209,210,209,211,211,211,210,208,211,212,215,213,206,213,203,199,170,215,214,207,194,213,150,212,188,133,130,16,102,86,100,139,118,98,147,105,56,46,73,87,118,92,52,99,56,55,91,117,97,62,92,44,66,106,92,82,98,113,101,87,102,102,106,86,111,48,81,82,118,106,84,96,54,85,144,104,109,54,87,118,189,174,114,160,125,120,83,233,227,193,168,87,167,203,226,228,159,158,78,221,215,188,156,89,174,41,29,177,170,128,105,204,209,187,175,133,159,181,217,208,170,121,105,218,204,185,167,147,180,194,201,202,179,136,150,197,197,179,173,163,210,198,206,172,161,128,162,210,192,176,64,89,58,143,193,157,145,154,199,207,214,175,130,163,176,195,208,112,130,119,122,185,193,157,131,158,142,156,233,207,190,57,110,91,191,56,102,51,118,55,63,92,108,167,185,215,109,82,83,79,122,40,179,126,53,77,124,145,70,157,75,125,
139,144,85,71,91,92,93,94,95,94,97,97,100,103,101,99,153,55,88,157,98,56,90,93,101,99,99,95,96,92,87,137,70,10,11,11,11,23,23,203,206,207,208,209,210,210,212,212,212,212,215,183,213,183,200,213,197,207,204,191,203,214,161,153,203,200,191,177,180,200,141,36,142,112,180,196,124,92,81,142,126,197,204,153,100,69,157,126,197,204,175,113,82,127,64,192,199,190,160,112,134,103,70,152,193,190,125,111,62,199,201,190,183,141,91,77,176,200,185,185,141,104,59,184,202,187,202,127,86,134,130,150,128,109,111,54,128,121,134,137,119,105,40,65,147,187,183,173,145,84,140,167,179,167,150,116,75,54,112,122,114,91,98,72,102,130,128,115,70,79,100,122,109,91,116,104,114,149,117,92,96,140,144,125,111,71,124,141,185,182,137,160,157,216,210,188,92,100,165,172,103,75,160,173,198,225,147,191,219,143,140,143,113,63,139,156,161,134,206,187,147,124,119,62,169,102,163,164,88,133,121,85,40,76,66,78,150,179,126,157,182,73,82,58,98,144,161,91,60,36,189,128,158,124,92,135,
142,146,85,88,92,91,96,93,94,94,99,99,99,103,102,99,152,52,89,157,99,49,90,91,103,97,97,95,97,93,88,142,119,10,11,11,11,12,65,206,205,207,208,209,210,211,210,213,213,213,212,214,182,196,179,213,215,214,215,210,213,192,212,154,152,175,183,209,174,187,28,162,117,168,91,118,56,59,103,157,162,151,102,102,62,76,77,159,150,113,119,83,58,57,150,165,144,127,101,87,81,71,91,135,165,120,94,76,127,175,172,172,110,92,87,69,106,156,155,148,120,107,79,132,145,118,136,117,85,62,165,144,139,112,102,98,72,184,200,174,169,154,115,99,178,174,202,201,166,126,143,167,164,221,206,177,127,139,173,170,203,201,173,132,113,191,218,204,198,154,125,123,207,199,189,166,142,188,199,211,202,180,137,148,216,209,196,178,138,201,205,204,185,159,138,182,174,102,104,142,111,174,192,114,223,220,193,172,141,124,112,195,107,148,170,157,150,85,142,142,100,161,95,143,144,105,128,110,144,79,121,50,41,101,87,58,93,75,162,124,165,110,95,89,65,117,127,63,47,172,113,78,94,108,185,81,
147,149,88,93,92,94,98,93,94,95,101,98,100,100,102,101,153,50,88,156,98,46,89,92,101,96,97,96,94,95,90,116,129,18,11,12,12,11,28,178,203,207,209,210,211,212,212,213,214,214,214,204,184,195,191,176,199,187,210,167,194,206,215,199,108,197,179,170,180,186,8,151,130,39,139,95,200,203,163,117,86,136,95,203,192,181,176,129,99,104,203,140,194,191,166,117,94,146,72,211,185,198,173,163,102,58,187,156,187,198,163,142,122,94,61,205,191,190,199,159,87,64,200,145,197,217,187,135,95,129,93,212,212,175,170,148,125,67,208,207,200,199,166,105,79,180,199,206,203,175,100,86,148,196,220,208,188,172,136,83,136,192,196,148,142,115,87,125,196,185,178,147,99,78,160,186,158,138,104,105,114,159,159,139,147,116,123,102,95,85,66,132,155,184,201,140,137,58,96,126,107,162,142,127,216,156,150,204,140,123,113,131,141,139,153,125,163,82,117,61,156,112,137,104,155,46,94,150,64,97,84,102,57,55,43,58,80,98,49,200,93,167,92,56,87,68,79,41,82,85,53,140,106,58,117,90,
139,127,89,93,94,96,97,94,95,94,102,98,100,101,103,102,154,41,87,155,97,45,90,92,101,97,97,97,95,94,90,86,136,80,9,10,10,9,18,34,207,208,209,211,212,213,213,214,215,215,216,217,213,216,205,193,143,189,205,160,191,217,209,193,200,165,182,142,188,120,138,92,57,38,92,132,127,124,98,115,57,70,192,199,175,164,93,78,66,82,115,184,192,165,127,97,76,55,152,197,196,143,155,104,81,127,97,201,215,178,159,119,72,58,143,116,184,199,159,132,117,84,84,74,111,130,155,123,118,117,54,69,113,128,132,97,78,63,101,93,93,89,81,104,55,91,77,140,136,130,112,103,113,68,182,164,157,182,147,130,130,158,186,214,212,183,161,136,173,134,217,208,189,164,153,160,179,216,214,202,182,172,170,162,216,216,194,172,160,208,188,197,195,175,146,172,205,171,112,132,188,145,192,159,165,125,153,168,141,166,99,104,121,196,206,163,190,113,111,57,73,124,32,48,99,56,93,94,189,98,86,82,35,109,87,85,78,135,160,143,115,177,166,107,88,70,87,104,62,50,171,172,86,62,188,190,
87,132,92,84,85,91,97,97,95,95,101,99,98,100,101,99,152,46,85,155,95,41,90,89,100,100,98,96,96,93,90,86,141,122,11,13,12,12,11,59,206,208,209,211,214,214,216,212,214,215,217,208,214,207,210,216,212,200,200,84,199,198,209,199,200,157,200,118,165,21,65,179,173,185,171,139,71,58,181,131,195,203,178,131,124,64,45,187,150,190,193,153,125,139,91,68,211,198,183,197,151,93,140,119,125,213,211,188,181,134,97,121,147,103,206,218,195,194,181,107,93,121,78,212,206,181,208,145,111,125,120,112,215,201,192,190,144,110,131,156,136,201,207,179,144,118,83,111,209,209,188,193,137,121,106,172,173,213,208,160,130,123,167,157,214,215,175,152,139,135,99,210,205,173,189,170,83,65,181,202,194,190,165,93,72,140,185,172,150,98,83,59,52,88,89,89,102,83,102,94,95,184,92,181,160,132,164,177,177,109,137,99,184,73,89,100,105,77,193,31,104,63,135,71,178,105,71,113,110,121,121,119,40,105,51,27,43,155,99,47,92,89,93,101,51,247,131,132,99,75,67,65,67,109,161,114,
45,79,69,74,84,100,94,95,97,98,100,99,99,100,101,99,151,50,80,153,93,34,87,89,98,102,98,97,98,94,91,87,122,126,17,14,12,15,21,43,195,209,210,212,214,214,207,196,199,217,211,211,208,217,217,219,217,219,216,205,216,206,153,202,203,178,75,192,146,42,197,102,92,42,77,78,158,114,83,110,85,83,39,55,48,52,36,42,30,21,12,7,12,11,16,17,22,10,13,10,10,12,11,12,9,14,11,12,15,10,16,14,13,12,13,11,11,20,14,12,15,32,29,47,49,63,42,23,58,37,65,71,86,81,98,83,61,56,31,77,99,128,156,103,126,71,115,83,178,182,208,197,156,120,93,109,75,198,199,183,180,149,106,78,157,169,213,206,181,165,154,128,99,198,209,201,189,170,126,140,177,192,212,198,170,108,120,210,196,196,187,170,128,116,192,213,193,177,102,105,120,173,195,184,161,112,207,138,194,121,190,47,136,66,104,161,150,211,32,18,30,30,197,171,85,67,73,125,150,105,155,156,72,105,41,70,77,61,57,79,43,69,47,30,52,145,211,150,118,67,202,127,51,88,57,152,
22,45,34,73,73,90,48,97,70,99,99,97,99,101,99,99,154,48,77,153,94,37,86,89,97,101,97,95,96,95,91,88,83,130,23,21,21,22,20,28,38,211,211,214,213,211,189,211,193,213,220,218,216,212,220,197,220,218,215,194,212,198,128,168,154,188,93,173,151,29,18,21,23,26,26,18,19,19,19,21,23,18,20,20,20,20,20,21,21,22,21,22,20,21,20,20,20,17,18,20,19,21,19,21,19,19,20,20,19,19,19,18,19,19,21,20,22,22,23,22,23,23,24,23,25,24,24,24,22,23,24,22,23,20,24,19,21,21,20,20,21,19,23,24,23,23,21,20,23,18,21,22,22,26,25,23,22,25,25,22,22,22,24,21,22,23,22,20,19,19,21,22,21,21,22,24,24,25,28,26,27,22,31,27,27,27,28,27,27,29,32,44,48,56,53,73,116,135,168,96,126,172,169,149,177,217,221,226,167,189,117,244,141,52,20,59,43,90,39,32,27,149,131,73,47,163,82,114,79,69,64,81,111,185,33,87,96,134,132,93,46,57,88,85,109,103,189,44,190,69,106,189,133,165,113,57,
21,13,26,49,66,30,41,78,56,94,100,99,98,99,99,91,148,49,69,155,95,33,84,83,98,97,97,93,95,93,91,89,87,140,20,18,19,21,30,10,49,208,212,214,206,214,213,188,188,208,209,212,219,215,220,214,219,221,206,201,213,216,168,217,105,173,203,177,159,65,124,193,84,160,200,86,172,98,93,93,17,85,60,42,49,50,49,51,51,51,47,55,52,54,54,54,54,53,56,57,56,64,54,59,57,57,59,58,59,59,60,61,61,55,58,63,62,65,68,71,51,77,79,81,84,86,88,50,88,95,99,98,99,101,103,82,106,110,111,113,113,45,111,112,113,114,112,114,50,112,112,111,110,111,114,65,111,113,112,110,110,111,110,27,106,109,109,110,109,109,99,40,98,94,87,74,72,65,26,53,48,44,39,34,30,24,23,20,20,23,20,23,26,22,24,19,23,18,18,22,118,176,147,134,165,127,124,141,87,100,188,96,43,51,72,63,99,68,41,42,32,130,191,75,65,174,104,141,125,45,109,118,167,86,107,72,32,86,53,66,87,72,49,104,60,44,59,63,90,99,45,164,131,109,114,79,
43,20,16,43,64,34,95,38,73,91,101,98,99,101,99,92,154,149,146,149,90,34,77,80,98,96,97,96,94,93,90,90,87,110,94,18,9,7,9,8,55,204,213,210,207,214,206,186,206,173,189,211,183,190,199,197,211,189,199,189,190,221,217,87,181,99,202,151,169,180,154,185,198,165,196,152,198,98,98,97,29,85,57,45,49,49,50,51,52,50,51,53,54,54,54,53,54,54,54,55,54,56,54,54,55,55,55,54,55,54,55,56,55,54,56,55,56,56,57,57,56,57,56,55,54,56,56,56,57,56,56,57,57,56,56,56,57,57,57,56,56,56,55,55,54,54,54,58,57,54,57,58,57,56,57,57,56,57,57,57,58,57,58,59,58,56,57,58,59,58,58,59,59,59,58,57,58,57,59,58,57,58,57,56,55,54,76,92,91,89,39,56,165,36,202,176,193,150,127,20,207,205,182,206,97,102,179,124,170,107,29,28,31,60,58,47,41,49,117,34,69,45,153,104,42,186,134,102,122,33,30,56,124,103,53,55,54,25,96,61,43,63,40,51,58,51,154,74,171,118,94,62,63,114,200,139,
77,10,12,21,16,34,63,48,94,96,100,98,97,98,98,90,130,148,145,153,97,153,135,86,96,98,95,95,93,94,92,90,89,82,123,12,6,9,9,10,21,40,212,217,201,203,211,183,218,222,219,213,202,197,212,202,201,212,209,216,171,208,212,155,149,118,156,71,150,165,211,207,174,141,197,187,197,75,77,76,54,18,49,46,49,51,51,53,52,52,54,54,54,55,55,55,54,56,56,56,56,57,57,57,55,57,56,57,56,56,55,56,57,57,59,57,57,57,57,56,56,56,59,57,57,57,58,58,57,58,57,57,57,57,59,58,58,58,59,57,55,57,58,59,57,58,57,56,56,56,56,55,56,61,59,57,57,57,56,55,57,58,57,57,55,55,56,57,57,57,56,55,55,54,56,56,54,54,55,56,54,53,53,52,52,51,95,90,90,86,51,53,186,40,125,130,147,97,142,136,208,193,162,129,179,83,112,91,26,51,72,16,35,105,151,37,40,26,67,45,56,139,138,80,85,49,155,212,31,82,34,80,39,85,51,37,65,28,108,84,48,46,49,33,150,30,101,60,86,98,131,153,88,148,173,93,
71,9,13,15,30,12,12,66,95,95,100,98,97,99,97,98,92,91,86,114,96,152,146,150,134,98,96,95,96,94,92,88,89,84,129,6,9,10,11,10,12,35,213,216,215,215,205,205,220,205,212,219,222,207,194,218,196,205,129,198,173,221,178,221,103,81,219,68,151,202,217,90,202,165,104,177,187,83,61,55,52,44,40,45,50,53,53,56,55,56,56,57,57,58,58,58,58,58,59,57,60,61,61,61,59,59,60,60,59,58,59,57,59,59,60,60,59,58,59,60,59,59,59,59,59,59,59,60,61,60,61,60,61,61,61,61,60,60,61,59,60,61,61,61,59,61,61,61,61,61,59,60,60,58,60,60,61,60,60,59,60,59,59,58,59,59,59,58,58,58,59,58,58,58,57,58,58,57,57,58,57,56,56,56,55,52,67,65,61,59,20,60,191,69,107,156,142,134,170,148,152,173,164,99,130,133,138,59,56,86,174,42,33,46,44,29,61,99,38,67,53,93,61,51,76,53,101,112,35,56,63,53,45,41,110,73,34,50,44,40,59,45,195,70,62,47,57,73,105,81,114,115,92,76,132,70,
66,6,5,8,44,13,20,35,96,97,96,98,98,98,98,98,94,93,94,90,89,84,83,146,126,96,95,95,95,94,92,89,91,85,137,8,22,11,12,11,9,54,188,203,195,193,213,221,223,214,198,156,195,220,207,213,193,207,202,151,128,102,214,212,154,127,195,173,195,214,176,123,181,189,73,206,160,158,77,59,56,55,27,45,55,57,58,60,59,58,61,62,62,62,62,62,62,62,62,62,63,64,65,65,62,63,63,63,64,63,63,64,64,65,64,65,62,64,63,63,63,62,62,64,63,64,64,65,64,66,63,64,63,64,63,64,64,64,64,64,62,64,64,67,64,63,64,63,64,64,64,64,65,63,62,63,65,65,65,64,64,64,64,65,64,64,64,63,61,63,63,62,61,61,62,62,61,62,61,61,60,60,59,60,58,58,52,53,46,30,26,56,171,172,167,152,171,182,196,95,182,154,100,163,37,107,37,51,20,140,35,88,69,65,122,100,94,86,56,87,37,52,23,29,57,60,91,48,143,66,33,101,45,30,108,51,159,107,65,48,52,60,195,50,98,47,131,109,47,88,110,57,71,73,96,57,
20,6,4,9,6,18,30,81,94,95,98,97,97,98,96,99,97,94,96,94,95,94,94,90,95,96,97,94,95,92,91,88,88,85,140,15,21,23,14,18,20,15,202,191,182,196,200,220,220,187,224,204,223,211,217,216,208,224,219,172,169,212,159,195,138,171,217,183,215,203,195,101,202,149,137,207,150,158,154,74,56,52,9,43,59,61,61,63,64,61,63,63,64,65,65,65,64,65,65,65,65,68,66,68,65,65,66,66,67,67,67,66,66,66,66,67,67,67,66,67,66,67,66,66,66,68,67,67,67,67,67,68,68,66,66,66,68,69,67,68,67,67,67,66,67,67,66,67,67,67,67,68,67,69,65,66,66,67,67,68,66,68,67,69,67,68,66,66,67,65,66,67,65,65,65,64,64,64,65,64,63,63,63,63,62,60,59,56,42,14,55,58,100,185,201,181,156,141,144,103,126,193,188,176,35,107,47,107,62,100,63,72,21,36,55,13,94,67,22,52,173,129,37,36,102,56,74,129,130,52,36,55,145,43,55,92,87,74,45,77,84,82,162,32,37,46,168,106,86,78,160,111,43,121,188,82,
51,14,4,8,8,7,24,52,84,101,98,98,97,97,98,98,97,97,97,97,98,96,96,92,98,96,95,95,94,91,90,90,90,85,138,213,216,190,115,214,190,165,208,165,212,195,221,203,219,217,214,212,216,225,208,199,198,216,202,197,165,146,137,187,206,79,186,193,91,190,159,180,135,160,181,205,140,157,159,156,73,58,13,46,61,64,65,66,68,69,66,66,66,66,68,67,67,67,67,68,68,71,73,70,67,69,69,68,69,69,68,69,71,69,68,70,69,69,69,69,69,69,70,69,69,69,70,69,68,70,70,71,70,71,70,71,71,72,70,71,70,71,72,70,72,71,70,70,69,70,69,70,68,72,70,70,70,70,70,69,69,69,70,70,70,69,69,69,69,70,70,69,68,68,68,67,67,68,67,68,67,66,65,65,64,64,63,57,23,22,57,62,43,92,180,183,161,159,172,149,140,225,177,156,101,121,72,41,37,124,44,31,96,31,17,23,20,94,73,54,53,55,57,49,48,115,67,96,32,42,75,49,27,145,46,109,79,72,180,67,159,60,72,39,51,108,131,113,50,55,139,87,43,93,167,138,
35,8,4,7,10,7,23,65,90,97,95,97,97,98,98,97,98,97,96,97,97,97,98,95,97,96,94,95,92,90,88,90,88,83,139,224,215,218,162,212,190,209,208,139,211,212,223,193,220,208,210,140,199,223,215,214,223,144,210,195,160,157,141,158,191,210,170,156,97,192,173,101,220,167,161,99,175,163,160,157,160,65,12,48,64,66,68,69,70,70,71,70,68,70,70,69,70,70,70,70,70,72,73,74,69,69,71,71,70,69,70,71,72,71,71,71,73,71,71,72,72,72,73,74,74,73,73,71,73,73,74,73,73,72,73,73,74,74,75,73,73,74,74,75,74,73,74,74,72,72,72,73,73,73,75,74,74,73,73,73,73,73,74,72,73,72,72,72,71,72,72,72,72,73,72,72,72,71,71,71,71,69,69,68,68,67,66,60,16,45,60,64,134,53,131,139,176,142,172,184,194,127,131,176,130,134,152,27,79,123,35,28,19,29,25,118,36,20,44,77,31,123,46,48,185,64,53,70,131,42,65,40,37,111,38,44,130,34,178,170,181,89,118,31,127,130,184,118,66,56,68,103,110,87,123,60,
9,6,1,8,7,15,47,37,78,96,100,96,97,97,97,96,98,97,95,96,96,98,94,97,97,95,93,93,93,91,88,89,86,84,142,190,223,215,178,181,204,211,205,213,216,160,207,184,225,223,193,213,195,214,168,218,194,178,223,217,206,182,171,226,226,166,114,137,177,175,158,83,197,198,226,168,211,162,161,161,159,161,16,50,65,69,71,70,71,72,74,71,72,72,71,71,73,73,72,72,72,72,74,74,71,71,73,73,72,74,71,72,74,73,74,74,75,75,75,75,76,75,76,75,76,76,76,76,74,77,76,76,76,75,75,75,77,77,76,76,76,76,77,78,76,78,76,77,76,76,76,76,75,77,77,77,76,76,76,75,76,77,76,76,75,75,76,75,72,73,73,74,74,74,75,76,76,75,76,74,73,74,73,71,73,70,70,63,18,46,64,67,134,133,68,135,113,155,156,184,150,125,174,128,127,146,97,124,152,42,35,50,24,90,31,52,95,27,43,90,36,139,43,87,58,61,111,40,42,52,24,52,32,47,63,39,87,131,66,216,120,60,53,51,59,79,125,60,39,76,112,35,70,105,152,61,
5,4,1,16,3,9,7,32,74,72,99,96,96,97,97,96,97,96,93,95,96,96,96,95,97,93,95,92,91,92,88,87,89,85,142,148,173,193,178,154,205,194,199,185,206,213,228,220,199,206,117,203,166,190,225,148,215,199,166,201,203,200,167,144,200,203,112,214,183,194,133,83,215,121,150,214,136,156,159,161,161,159,55,52,69,72,74,74,74,75,74,74,76,76,75,76,74,74,73,74,73,75,77,76,75,74,74,76,75,76,76,74,77,75,76,77,76,76,78,77,77,78,78,79,79,78,77,77,78,75,76,77,77,76,76,77,78,77,79,78,78,79,79,78,78,79,78,79,76,79,77,77,78,76,77,77,77,78,76,77,78,79,79,78,75,76,77,76,75,75,75,73,73,73,76,76,78,76,76,76,76,76,74,75,74,72,72,67,20,48,67,69,147,135,140,168,121,177,75,157,160,201,72,143,110,150,150,38,79,26,35,16,29,55,25,32,45,54,19,26,39,58,65,93,64,69,47,71,33,21,32,56,89,30,52,38,63,145,106,76,76,59,88,68,80,83,77,156,88,64,49,76,47,87,88,82,
2,1,8,9,5,4,10,101,28,56,97,94,98,98,98,97,97,97,94,96,94,95,95,94,96,92,92,91,90,92,91,91,87,86,139,138,183,187,194,167,195,173,153,163,188,191,187,221,179,145,203,210,189,174,227,222,201,205,168,204,159,126,153,137,202,167,207,178,200,110,163,89,136,135,182,118,158,167,165,177,160,162,71,54,70,72,76,76,77,78,77,75,77,76,76,78,76,73,73,76,75,75,75,77,75,78,76,78,78,77,77,75,78,78,77,78,79,79,80,79,78,79,79,80,79,79,79,79,77,76,77,78,77,76,76,76,77,79,80,80,80,80,80,80,79,79,81,81,79,80,80,78,78,77,77,77,77,79,79,77,80,80,81,80,79,80,80,77,76,77,75,77,77,77,78,79,77,76,76,78,79,76,79,77,76,76,73,70,22,49,70,72,127,146,101,140,101,165,80,190,118,109,20,126,55,62,45,149,59,22,25,39,25,59,30,106,21,20,29,39,28,135,56,39,89,188,50,75,42,30,19,59,88,47,39,26,64,49,75,52,60,82,110,67,80,177,60,103,120,54,72,35,43,124,118,35,
1,1,0,3,3,6,68,40,29,22,94,87,93,95,96,98,94,95,93,94,95,94,94,93,94,94,92,91,90,92,91,91,87,86,141,181,142,173,173,143,183,187,171,168,190,163,133,151,149,147,181,200,219,185,196,217,229,177,114,163,150,191,193,165,164,172,148,108,111,66,142,144,213,170,165,161,192,172,168,165,167,169,70,55,72,75,77,79,78,79,78,79,79,78,77,77,77,72,62,124,127,100,66,73,78,78,79,80,80,79,80,79,80,80,80,81,81,80,82,80,82,81,81,81,81,80,80,80,79,78,78,73,73,72,71,72,71,77,80,81,81,82,85,82,81,80,81,83,81,81,83,78,79,78,77,77,80,81,81,79,80,81,81,79,79,77,73,71,73,75,78,78,78,77,79,79,81,81,81,80,79,78,80,79,79,80,78,72,22,49,71,75,112,115,145,158,158,138,131,119,144,135,34,79,146,23,25,34,153,35,47,23,29,23,32,30,128,66,62,56,31,43,58,75,166,137,59,50,34,89,54,37,42,23,45,56,52,46,69,34,50,37,30,88,38,80,197,87,47,54,162,47,60,173,107,63,
1,0,3,1,2,3,32,23,19,53,63,77,92,96,97,95,95,94,92,94,95,94,94,92,94,92,93,91,90,89,89,90,88,85,141,148,118,167,191,163,197,189,178,162,190,185,130,136,135,161,128,113,214,169,210,156,197,214,167,121,145,156,211,173,179,156,179,98,195,90,168,119,187,229,160,184,200,144,162,163,162,165,80,57,74,77,80,79,79,80,81,80,80,79,79,76,141,142,140,141,142,138,140,141,119,72,81,80,82,81,81,81,80,81,82,83,82,82,83,82,83,82,82,83,83,82,80,81,77,80,76,146,142,144,146,146,148,146,81,79,84,83,85,85,85,82,84,84,82,82,84,80,79,72,68,72,79,82,82,84,81,83,84,80,73,83,145,138,140,141,146,76,73,76,80,81,81,81,80,80,80,80,82,81,80,79,78,74,23,51,71,76,118,112,123,156,149,142,137,48,93,48,92,131,147,35,60,81,154,18,49,24,31,38,23,58,38,25,13,56,43,173,95,158,121,76,80,37,53,31,62,33,22,29,61,44,49,152,51,28,53,42,50,67,64,109,211,69,71,57,40,51,49,118,87,86,
3,2,2,2,2,5,9,10,60,121,54,83,147,100,95,92,95,94,93,93,94,94,93,92,95,91,92,90,89,89,90,90,87,84,141,165,157,149,197,147,206,174,180,162,117,135,156,136,151,134,130,117,93,100,173,165,147,198,185,164,139,187,150,99,117,145,169,100,109,127,162,73,140,164,119,114,201,158,162,167,164,165,85,58,75,78,80,82,81,81,80,81,80,81,78,143,143,139,139,138,136,140,136,139,136,141,79,82,85,84,84,82,81,83,80,83,83,83,83,84,84,83,83,85,85,84,82,82,81,116,147,143,140,140,141,138,142,144,147,140,82,85,85,85,85,85,85,87,86,83,85,81,76,139,141,140,137,76,86,84,85,83,83,67,141,140,139,137,135,138,139,139,141,93,82,82,83,82,83,83,83,81,80,81,81,81,81,74,23,51,73,78,121,117,118,141,138,153,151,155,85,54,83,143,127,51,74,80,42,40,24,24,36,37,76,85,37,40,21,24,29,102,81,121,47,103,51,58,36,134,26,35,98,32,48,38,28,115,53,110,79,34,99,72,71,50,189,48,191,47,29,43,118,151,127,35,
1,1,1,1,1,2,16,10,10,36,117,133,148,102,96,92,93,94,92,94,93,92,93,92,94,90,90,91,88,89,89,88,86,83,141,154,162,174,138,153,156,165,179,133,162,161,142,171,141,168,166,123,100,133,132,115,134,113,171,119,136,104,136,140,75,155,91,81,84,101,146,81,202,205,123,198,194,155,167,170,159,170,85,58,75,79,80,178,82,81,79,82,82,81,80,143,140,118,28,16,10,23,37,131,136,142,89,81,85,86,84,84,83,85,85,82,83,83,84,84,85,84,85,84,85,86,83,83,82,147,142,134,54,19,14,22,65,139,146,146,78,85,86,86,86,87,87,89,86,87,84,82,134,44,16,23,94,134,83,85,84,83,80,145,140,137,128,105,90,130,137,137,141,147,70,83,85,84,84,84,82,83,83,84,83,81,81,76,19,47,73,78,121,121,117,132,118,194,91,81,56,54,89,34,39,133,23,93,43,63,32,115,20,25,26,124,23,37,93,75,38,34,47,122,40,133,54,38,47,153,28,34,78,114,34,42,67,158,111,34,47,30,39,56,51,52,152,22,208,173,37,58,185,159,57,25,
12,1,1,1,2,43,7,7,59,113,135,146,110,90,95,93,92,94,93,93,92,92,94,91,91,92,90,92,93,90,87,87,86,84,140,193,172,127,164,182,160,159,168,143,147,157,144,148,126,166,138,165,148,76,110,151,97,125,170,166,129,95,204,140,171,182,152,76,157,193,85,105,164,152,227,183,197,161,173,168,165,171,94,59,76,80,81,167,176,86,80,82,83,84,80,138,123,14,23,25,13,19,14,16,11,143,114,81,84,87,85,85,84,83,85,84,84,85,87,86,85,84,84,86,85,85,85,86,81,143,24,16,20,12,16,21,18,12,28,145,81,84,87,87,87,87,88,88,86,87,86,81,136,4,3,2,5,140,83,85,86,86,82,146,74,14,7,4,9,18,20,25,112,145,77,85,86,86,84,84,84,84,85,87,84,82,77,77,23,52,75,79,163,125,118,124,113,166,164,88,89,68,43,93,93,45,24,130,26,35,44,45,27,62,28,137,21,53,26,96,18,45,118,89,53,103,23,30,110,82,30,24,55,56,29,40,85,32,138,51,23,35,105,35,44,97,91,20,160,66,31,69,127,43,25,40,
4,1,0,1,1,29,28,24,18,18,17,58,76,50,58,91,92,93,93,93,91,91,93,91,91,90,145,133,94,131,88,88,86,80,138,200,133,174,188,166,167,183,154,110,160,171,156,170,192,165,118,134,100,141,70,86,61,72,97,101,140,177,159,161,169,198,149,116,110,159,75,148,189,95,185,220,178,173,173,178,165,172,75,60,75,79,84,185,183,176,83,81,83,84,81,141,125,13,28,24,15,19,21,11,12,144,113,83,85,86,85,85,85,84,85,85,86,86,85,87,84,87,87,87,86,88,85,85,82,144,17,10,7,9,15,8,11,20,13,145,81,86,88,86,86,87,87,89,88,86,87,84,135,1,2,2,8,139,85,87,86,84,79,143,38,3,3,3,13,18,19,13,41,143,78,85,86,87,85,85,84,86,85,87,85,85,83,76,24,53,76,80,127,162,138,140,178,167,111,167,59,98,116,160,69,20,19,41,33,27,23,53,47,58,50,78,39,58,23,30,12,25,40,49,71,25,48,24,119,78,42,100,60,44,23,145,38,34,79,32,47,82,71,160,33,48,65,42,49,91,90,54,22,45,53,142,
1,1,1,1,2,5,15,4,72,14,16,32,126,81,93,91,92,93,92,92,91,91,92,91,89,90,145,145,141,141,87,87,86,82,138,123,165,167,162,171,159,163,133,124,149,175,118,136,105,156,151,153,88,70,86,124,98,143,152,149,215,154,121,113,182,116,174,181,136,198,66,88,161,193,145,222,132,169,175,177,178,171,75,62,79,81,86,176,182,176,176,87,86,84,80,139,124,14,30,25,17,20,32,11,14,143,115,86,85,86,86,84,85,86,86,86,86,86,86,88,87,87,87,86,87,86,88,86,84,140,16,11,8,10,16,10,11,12,15,146,80,87,88,88,87,89,88,89,89,86,87,85,137,2,2,1,10,140,85,88,88,84,78,138,41,3,3,3,12,23,30,17,54,142,80,85,87,85,87,87,86,87,86,88,85,85,84,77,25,53,75,79,157,166,118,171,155,175,37,120,81,111,51,90,157,102,31,37,32,25,14,24,58,33,69,89,40,32,33,36,25,48,33,47,66,50,46,49,35,50,183,77,53,27,39,51,78,140,132,49,50,91,86,55,50,27,56,144,129,84,21,27,28,56,156,192,
0,1,2,2,31,22,4,1,3,9,8,48,87,92,93,89,91,91,91,94,91,90,90,91,90,90,140,135,141,141,87,87,83,84,132,190,173,182,95,154,171,191,163,172,161,152,161,135,85,103,98,171,154,159,169,76,147,133,134,116,130,152,164,155,93,115,137,138,167,134,40,132,102,92,99,168,141,174,182,170,169,172,89,63,79,81,88,180,177,179,177,166,88,85,83,140,116,18,34,24,17,31,14,12,15,143,115,84,87,87,85,88,86,87,87,85,86,86,85,88,87,89,87,88,87,88,86,88,83,140,14,13,8,10,16,10,15,27,15,146,79,87,88,89,89,89,88,89,88,85,87,85,136,2,1,1,9,136,85,89,86,84,81,138,40,3,3,2,13,21,19,14,56,141,81,84,87,88,89,87,86,88,86,86,85,85,83,79,25,54,79,81,48,183,154,147,142,177,119,191,83,108,77,55,126,87,13,11,19,27,10,33,39,41,72,155,41,36,67,60,23,36,13,57,52,19,84,66,36,75,83,46,96,38,50,110,149,146,156,80,56,79,79,203,66,44,57,75,85,25,27,41,39,156,186,155,
1,1,1,33,41,2,4,2,47,7,13,87,139,93,89,53,74,82,94,93,92,90,91,93,91,89,142,14,58,82,86,84,84,82,133,176,176,178,154,172,150,166,132,165,148,170,177,136,175,171,95,128,160,142,64,93,116,177,82,123,143,81,134,113,84,148,111,124,163,98,37,171,121,115,98,192,192,175,176,169,169,175,95,64,79,82,86,180,176,177,179,178,159,86,81,142,104,12,16,15,12,21,14,12,13,144,118,87,87,88,88,87,87,88,87,85,85,87,86,88,85,90,87,86,89,88,88,86,84,140,15,15,9,12,15,14,17,29,15,145,80,86,88,91,91,89,90,89,89,88,89,85,139,2,1,1,11,138,83,87,88,87,83,140,40,3,3,2,14,13,19,14,42,140,83,85,87,87,87,87,87,87,88,88,85,84,84,77,25,54,76,80,49,220,197,190,172,156,140,113,117,42,29,27,95,84,23,23,41,19,22,60,77,101,132,128,37,31,79,52,20,92,59,68,96,27,47,24,27,42,156,44,132,66,93,48,157,79,161,88,76,106,34,43,48,48,46,46,50,21,41,65,117,141,134,191,
1,1,5,5,1,1,15,6,31,27,19,87,143,91,76,30,74,91,94,92,93,91,90,93,92,89,139,19,71,88,86,84,81,83,129,152,161,154,174,194,160,168,151,146,136,137,101,134,104,138,98,88,122,135,120,150,84,99,60,94,111,127,94,136,80,92,55,93,86,61,49,98,149,183,76,78,162,173,172,170,175,176,88,65,78,83,86,183,174,180,179,176,177,156,83,142,100,14,18,19,12,16,15,10,11,145,118,86,88,86,89,88,88,87,86,85,88,86,89,90,88,89,89,88,88,87,87,88,83,142,15,12,15,18,15,20,20,21,14,146,78,84,88,91,90,88,89,89,89,88,88,85,138,2,1,0,9,138,87,89,88,88,81,138,41,3,2,2,13,21,18,16,50,144,81,87,87,87,86,88,85,87,88,86,85,83,84,77,26,52,76,82,35,234,189,200,201,129,205,155,46,24,48,157,63,48,21,17,25,20,112,33,36,122,107,112,50,31,85,113,39,40,43,31,48,113,19,27,19,54,204,55,180,214,200,84,54,136,38,147,17,21,42,50,35,148,67,39,45,65,69,54,74,223,157,176,
0,5,1,3,2,14,32,44,109,47,20,87,146,85,54,55,51,43,83,94,93,92,91,91,90,89,138,23,76,89,86,85,82,94,131,139,131,120,187,181,179,135,153,126,160,133,130,164,125,205,67,84,107,84,52,74,106,115,73,148,78,111,112,78,37,121,147,189,158,117,52,33,93,171,82,170,100,176,166,169,174,172,80,66,80,82,83,181,178,181,177,169,179,181,130,140,116,15,17,15,16,19,12,11,15,144,107,85,87,88,88,86,89,86,88,89,86,87,89,88,89,91,89,91,90,88,90,88,84,140,18,7,13,13,15,5,13,17,15,143,81,88,89,88,91,90,89,88,89,89,89,86,137,2,1,1,10,140,83,87,90,90,84,139,37,3,2,2,13,22,19,19,27,143,80,87,86,86,87,87,85,87,86,86,85,85,83,77,26,54,78,81,43,238,214,192,199,179,119,141,51,15,28,42,85,144,28,11,20,24,89,105,22,143,58,65,83,88,88,111,55,60,57,93,112,50,23,37,39,55,212,155,37,179,114,237,220,82,68,150,64,43,44,59,41,12,72,23,165,188,77,75,168,140,188,94,
0,6,5,41,50,22,47,96,147,25,20,91,142,74,45,13,51,46,84,69,92,91,91,90,91,89,137,23,78,92,84,84,84,94,129,124,138,144,153,138,151,137,125,155,152,172,149,151,97,108,62,118,91,104,102,51,58,88,65,69,40,48,41,87,73,133,137,136,143,157,128,140,74,77,127,123,104,171,169,171,183,173,79,67,79,82,85,176,179,184,180,174,180,183,170,154,118,17,37,21,14,16,9,12,13,143,101,86,87,89,87,86,86,87,87,89,88,90,90,87,89,89,90,90,89,90,89,88,82,140,19,6,13,13,16,6,10,11,17,140,81,91,91,87,90,91,91,89,89,89,88,88,133,0,0,0,8,140,88,90,89,88,86,138,42,2,0,0,14,19,13,13,28,145,81,84,87,87,88,86,88,87,87,85,86,85,84,77,27,53,79,82,20,237,218,182,197,198,227,153,49,25,61,89,65,19,17,14,13,71,37,50,38,155,38,84,55,27,74,122,77,36,32,36,129,61,36,61,29,49,136,179,111,214,199,148,71,31,72,114,37,37,60,66,45,19,77,155,150,115,148,78,89,178,116,86,
2,4,8,9,14,31,16,56,92,48,27,90,117,63,11,11,48,14,49,41,60,83,92,88,90,88,136,23,82,96,85,82,83,94,124,96,93,222,125,104,124,97,119,118,106,140,134,84,129,193,111,109,124,145,114,108,57,55,40,40,79,134,63,129,87,120,160,58,108,49,176,39,167,67,122,114,133,168,172,172,177,173,82,68,79,84,84,172,180,180,171,178,181,176,165,206,131,18,39,39,17,16,9,13,13,138,100,87,88,88,88,89,86,87,89,88,89,91,89,89,89,88,90,89,89,89,89,89,84,139,18,5,12,11,16,6,12,12,17,144,82,89,88,89,90,90,88,89,89,89,89,85,135,0,0,0,7,137,87,88,89,90,85,138,41,2,2,1,15,15,11,11,22,142,80,85,86,86,87,88,90,89,86,85,85,83,84,78,27,55,77,81,22,174,187,202,195,200,206,157,68,39,25,33,24,31,11,62,21,77,29,164,98,93,46,53,56,45,35,65,69,47,36,29,107,103,49,69,30,53,55,45,159,104,209,80,57,90,43,114,25,30,44,39,51,35,64,143,43,184,146,78,124,105,179,180,
4,48,22,31,23,11,68,69,121,52,24,90,121,26,14,10,68,37,35,71,59,82,91,87,89,87,136,17,80,102,81,80,80,98,120,116,156,141,112,132,103,79,179,145,130,140,155,150,136,194,106,114,91,77,95,78,44,64,64,49,67,148,111,126,137,93,78,99,93,100,158,29,77,35,76,108,124,168,171,175,172,173,91,69,82,85,89,177,180,177,177,176,183,175,173,205,144,17,44,40,16,16,9,16,12,141,98,89,89,90,90,88,86,89,88,87,87,89,89,87,90,90,90,90,88,89,89,88,84,135,17,4,13,12,16,7,13,15,16,138,81,88,89,90,90,90,89,90,89,90,89,85,128,11,10,11,14,133,86,87,90,91,86,139,40,1,2,1,15,15,13,10,43,141,79,89,86,87,90,89,89,89,88,87,86,86,84,77,27,54,79,80,35,249,189,194,186,123,229,150,34,82,25,43,31,21,24,97,37,35,73,150,87,106,71,57,40,28,42,32,69,19,17,35,58,110,94,45,27,108,213,173,127,162,190,209,55,61,39,71,59,58,62,26,66,51,190,178,118,68,74,67,82,93,113,193,
2,40,9,12,16,57,65,65,119,51,34,89,108,15,11,18,35,25,51,43,66,63,87,85,89,87,135,23,84,109,83,82,80,104,137,240,230,141,225,178,196,168,111,188,129,196,212,146,178,127,123,160,209,130,178,51,70,89,65,88,125,111,117,83,174,117,93,116,104,90,94,48,59,133,151,58,113,168,177,170,171,175,95,70,81,86,90,178,178,181,180,176,185,171,172,196,154,18,29,32,15,16,8,15,13,137,95,89,88,88,91,88,88,90,89,88,86,88,89,87,89,92,90,89,88,89,87,88,83,138,16,6,11,11,15,10,21,24,16,139,84,90,90,90,90,92,88,90,90,87,89,84,99,47,41,34,31,102,86,88,89,89,88,138,42,1,2,0,15,17,12,11,59,142,79,89,89,87,88,90,90,90,88,88,87,85,83,79,27,54,77,80,18,249,192,197,84,104,225,121,45,49,35,23,75,20,21,63,102,58,32,85,138,67,74,74,62,11,26,53,61,27,58,24,32,72,75,61,62,88,69,129,119,160,200,148,41,106,56,60,89,61,86,43,43,47,142,85,191,56,50,65,171,154,204,142,
1,8,4,8,20,44,30,36,105,53,25,57,94,18,5,31,32,21,28,22,66,87,89,85,88,87,133,24,85,112,81,80,78,105,132,223,200,233,110,201,196,131,62,145,156,182,118,120,192,131,67,146,104,116,162,106,69,95,132,110,102,114,76,182,68,96,98,104,56,75,102,62,89,135,80,115,118,164,177,168,173,181,86,71,83,87,93,179,180,181,179,178,178,158,170,203,138,21,29,25,15,18,12,15,14,140,93,88,90,90,86,89,88,90,88,89,89,91,90,85,90,90,90,90,90,88,88,88,87,138,16,7,11,11,16,11,11,18,16,144,86,90,91,91,90,92,92,91,92,90,90,88,146,142,148,147,144,147,82,89,91,91,87,139,42,1,1,1,14,18,12,9,68,141,83,89,89,89,89,90,87,85,86,88,88,86,85,79,28,54,78,81,22,252,197,192,84,79,40,146,78,27,27,42,62,20,26,19,113,27,37,75,133,85,31,37,175,26,17,33,43,16,40,20,61,68,59,95,65,71,69,134,91,170,177,220,156,229,59,92,51,57,30,41,43,68,171,119,95,103,108,48,121,144,65,88,
3,10,3,9,8,20,32,28,74,50,25,34,35,7,5,2,3,19,30,54,76,84,88,85,88,84,132,21,84,119,80,80,78,105,125,121,126,120,133,158,117,110,76,120,73,87,132,122,121,96,94,118,89,111,95,114,46,62,137,128,118,71,116,123,126,117,74,104,169,155,93,75,122,79,75,135,151,167,171,172,176,172,83,73,83,86,96,180,179,183,174,176,177,167,180,206,143,21,35,29,14,17,13,13,14,141,93,89,91,90,90,89,90,90,91,88,90,90,89,89,91,93,89,91,90,90,90,87,85,137,16,7,9,12,15,11,9,11,19,143,85,91,93,92,93,92,93,90,91,90,92,90,119,138,145,149,146,146,87,91,91,90,88,139,40,1,2,3,14,17,15,13,65,145,82,90,88,89,91,90,91,90,87,87,87,87,86,80,28,55,77,81,59,252,228,205,105,153,90,164,52,18,46,79,35,17,136,61,119,28,93,138,90,32,48,30,95,46,45,69,43,36,14,21,84,126,47,74,75,89,54,112,64,85,118,191,152,239,142,68,45,44,22,25,31,51,103,140,165,154,90,84,173,140,113,153,
4,29,3,8,11,8,12,50,100,41,18,9,11,15,2,1,7,34,9,76,86,87,88,86,87,84,132,22,85,122,79,79,78,109,132,161,151,245,98,176,233,226,180,118,113,208,236,206,210,141,96,137,129,162,211,96,112,105,101,87,79,133,176,221,170,164,105,120,88,50,124,57,131,54,49,73,104,165,168,172,178,183,79,74,84,87,94,184,181,181,177,175,172,170,176,201,145,15,16,16,17,20,19,16,12,143,85,90,92,91,90,92,89,90,91,89,91,90,90,91,91,92,91,92,91,91,91,90,86,138,15,9,11,15,15,13,11,11,19,142,84,91,94,92,92,93,94,91,93,92,94,90,93,91,93,92,93,90,91,92,91,92,88,139,39,1,0,5,14,22,13,11,75,145,82,90,90,90,90,91,90,88,90,87,88,88,86,78,28,55,77,82,194,187,188,185,137,189,197,194,37,20,27,72,73,47,81,88,48,78,39,94,121,24,66,150,76,26,65,54,49,26,33,15,132,92,30,100,78,45,38,39,58,37,126,153,56,124,48,35,44,63,34,29,39,45,117,202,211,207,104,74,167,124,84,117,
3,4,2,1,21,10,18,49,92,22,5,19,3,5,2,3,7,23,64,82,87,86,86,84,85,84,133,23,85,124,81,79,78,111,123,183,134,233,222,148,192,221,190,136,125,206,221,168,141,145,64,78,65,98,95,178,129,221,64,126,167,168,193,149,167,89,170,66,56,62,136,85,122,78,49,72,117,165,179,178,173,181,80,73,85,87,96,185,179,177,178,173,174,170,176,201,143,26,25,16,13,24,21,14,11,146,87,89,92,91,89,92,90,91,91,92,91,92,91,90,90,91,92,90,92,93,91,89,86,139,15,14,18,16,16,18,17,16,21,140,86,89,91,91,92,94,93,90,93,92,94,93,94,93,96,95,97,96,93,92,92,92,88,140,36,1,6,6,15,18,17,19,85,147,81,90,91,91,91,90,88,87,90,88,86,87,85,80,28,55,78,82,142,147,142,140,143,180,156,186,61,54,40,81,48,21,29,91,41,17,42,71,21,21,38,150,74,58,71,58,75,36,26,39,107,115,46,137,123,21,36,49,160,42,86,136,86,79,73,53,106,69,56,38,26,47,67,160,125,101,153,75,115,63,129,131,
2,34,0,4,4,1,23,63,55,23,1,10,3,6,3,7,17,24,49,89,88,86,86,84,87,83,132,22,84,124,79,78,77,112,140,186,188,223,240,175,178,243,212,200,152,184,222,147,231,199,179,173,164,149,229,149,162,47,188,229,172,184,95,214,180,90,68,83,140,62,38,158,49,167,59,55,41,162,174,181,178,183,82,74,83,85,97,181,178,176,176,171,177,178,174,206,133,24,34,33,15,18,14,15,15,146,84,91,93,92,90,92,91,92,93,91,93,94,93,92,94,92,93,91,93,93,91,89,88,142,16,16,15,13,16,9,9,10,21,142,86,92,93,92,93,93,94,93,92,93,91,95,94,96,93,95,97,94,94,93,93,93,89,141,39,1,7,4,14,20,15,14,87,146,81,89,92,92,93,90,88,88,88,88,87,87,85,81,29,53,78,81,202,199,197,197,199,117,205,195,16,77,91,112,47,40,23,26,160,21,87,72,22,20,15,164,95,142,68,42,51,73,11,46,147,119,43,183,136,19,27,56,70,101,36,177,215,112,85,107,66,87,21,28,32,49,166,75,147,170,169,125,86,71,105,78,
3,5,6,5,8,4,4,61,26,12,0,6,3,2,2,7,11,33,88,87,87,86,87,83,86,83,132,17,84,124,79,78,76,112,129,84,232,195,150,158,197,91,197,166,140,182,161,198,163,179,118,157,144,129,217,191,60,180,82,168,191,185,150,57,111,206,87,68,110,91,86,61,47,116,96,29,42,163,181,176,179,182,79,73,84,85,105,179,180,181,179,179,176,176,178,206,117,28,37,15,15,19,15,17,22,159,84,90,93,90,92,91,91,92,92,92,93,94,95,94,93,94,95,93,93,91,92,89,89,138,17,14,12,17,17,6,6,6,23,142,88,91,93,94,96,94,92,91,93,93,92,94,93,90,92,95,96,95,93,92,92,93,89,140,43,2,9,5,17,17,16,14,92,144,82,88,92,90,89,90,90,88,90,89,87,85,85,80,30,51,77,83,210,202,200,198,188,221,202,102,42,33,115,57,33,52,16,60,61,31,76,52,52,83,28,115,114,121,89,45,82,105,115,118,196,40,148,133,147,24,61,134,150,173,163,196,187,117,87,105,175,49,15,43,48,26,32,59,93,164,164,75,84,92,119,76,
3,8,4,5,3,5,9,50,6,10,1,3,2,2,7,14,27,71,73,86,87,86,85,83,85,82,132,21,84,125,78,77,75,111,146,139,194,99,179,135,159,176,223,117,218,164,193,189,220,239,144,185,194,150,238,116,222,162,223,229,215,151,112,131,142,78,128,62,54,67,30,75,35,103,99,34,49,171,184,167,175,174,84,75,83,86,107,179,181,182,181,179,178,172,178,203,96,31,34,16,15,20,18,18,28,223,84,92,93,95,94,92,92,93,94,95,96,94,95,94,93,92,94,94,89,91,91,85,87,139,19,18,18,16,17,4,7,8,23,143,88,94,96,95,95,94,95,95,94,93,95,94,93,92,95,95,96,96,93,91,92,93,89,143,41,2,9,6,15,18,20,17,87,144,83,90,92,91,90,91,91,89,88,91,90,86,84,80,45,54,76,83,229,233,233,238,234,231,228,213,30,92,111,35,110,28,15,98,22,61,152,21,71,114,71,122,82,106,71,89,63,181,209,201,210,63,43,141,131,66,38,117,147,151,153,198,154,115,68,116,73,153,24,38,41,29,31,92,157,146,190,157,76,90,84,64,
4,3,3,4,17,10,36,69,11,7,1,2,1,1,9,20,27,47,87,86,86,86,85,82,84,80,130,20,85,124,77,76,76,110,160,192,242,148,237,191,240,52,177,155,177,199,215,205,225,158,216,146,211,194,169,212,139,229,149,183,173,69,150,110,132,125,87,88,136,127,76,80,50,41,84,74,63,165,182,175,174,172,90,75,85,86,119,178,180,183,186,178,174,168,171,206,89,28,23,14,17,28,21,19,31,221,97,160,145,119,110,99,94,94,95,94,92,94,94,93,95,95,93,95,92,93,93,92,91,136,19,8,12,14,18,6,9,12,22,142,89,95,95,96,95,95,96,95,94,94,96,94,95,95,96,96,98,98,94,93,93,94,91,140,39,3,10,7,16,21,20,17,84,148,91,92,92,93,93,93,91,90,91,92,91,86,88,84,81,53,77,83,158,157,158,159,161,159,163,163,95,108,141,42,85,24,10,76,22,130,129,37,65,19,56,95,95,115,45,68,24,172,184,184,187,128,33,81,66,119,39,124,150,189,154,190,164,80,69,86,87,58,37,39,44,42,20,95,77,157,126,91,139,99,68,67,
5,0,3,3,6,20,57,70,20,2,1,7,1,2,2,12,24,52,89,86,86,85,86,83,84,81,130,19,85,121,76,75,73,111,133,241,152,239,229,164,241,105,241,125,214,29,103,213,170,205,147,220,207,137,232,173,237,147,168,137,160,145,188,72,66,94,123,160,95,67,47,40,30,164,90,83,50,177,184,173,176,178,82,75,84,89,146,182,184,185,182,183,178,170,171,196,89,29,18,14,17,26,25,19,31,225,94,167,185,178,174,167,150,138,121,115,105,100,95,95,96,96,98,96,96,100,102,102,104,171,22,5,3,5,18,8,7,18,24,140,89,97,95,96,96,95,96,94,92,93,96,93,94,96,97,99,99,99,96,95,94,96,94,163,48,2,11,7,19,25,25,17,91,204,100,119,112,122,125,118,115,120,113,113,105,105,99,91,102,54,79,84,131,127,125,127,126,126,121,124,100,102,108,62,84,35,42,94,38,33,51,36,70,83,78,61,117,97,74,74,53,112,119,121,123,96,28,119,62,28,56,59,121,184,154,186,169,94,85,42,64,85,58,80,83,99,48,65,170,70,135,96,86,57,110,101,
4,11,3,6,5,5,19,61,11,3,2,2,24,2,5,67,59,86,87,86,85,85,84,83,82,79,127,18,84,122,77,74,74,114,174,208,175,231,237,222,168,227,160,234,151,142,92,134,227,126,231,162,190,104,160,239,203,148,142,99,185,93,79,50,79,137,75,43,81,95,87,51,23,184,62,70,30,181,172,172,179,179,85,77,85,91,146,183,182,182,180,180,179,178,178,208,76,27,10,21,17,48,46,22,34,227,95,173,183,176,179,182,177,180,180,179,170,158,160,154,147,145,149,152,148,158,159,157,162,204,21,10,5,5,18,8,8,17,26,192,91,111,106,106,105,106,102,103,107,106,104,101,100,101,104,105,104,110,116,122,122,128,140,204,56,3,10,7,19,19,28,20,87,227,99,165,164,167,167,171,171,166,169,166,167,153,162,156,129,56,79,85,156,172,167,175,173,175,168,172,123,83,47,72,119,148,56,135,104,34,156,159,89,152,145,162,151,41,26,109,162,164,162,178,118,52,18,23,83,12,56,130,116,127,138,156,108,143,90,43,104,164,52,42,83,45,20,109,63,42,94,128,137,73,80,64,
3,2,5,2,3,10,9,38,5,4,1,4,18,1,12,60,84,84,86,86,86,84,83,82,83,78,127,18,83,121,75,75,73,114,103,50,51,55,51,129,52,53,181,76,35,20,24,48,26,34,69,44,61,98,136,129,112,106,131,69,138,123,61,59,47,49,30,62,72,80,57,115,47,200,49,49,29,185,176,164,181,183,68,76,87,93,145,185,182,180,183,182,181,183,189,212,77,32,8,14,14,61,36,25,29,226,101,177,186,181,182,184,183,186,185,189,184,186,183,187,187,185,186,186,180,181,184,183,186,209,19,24,9,7,16,12,33,19,25,215,95,171,160,158,161,165,159,153,158,163,162,161,156,158,162,165,162,165,163,170,172,171,181,209,60,5,9,7,19,40,67,37,90,217,109,179,181,184,181,182,184,179,182,179,179,180,180,178,152,56,81,86,169,209,185,181,172,162,225,215,98,54,70,46,58,80,107,55,33,22,32,99,106,124,121,109,85,41,25,19,124,124,121,120,68,28,42,30,18,55,69,64,26,62,152,130,80,68,84,126,181,122,65,35,24,29,5,97,74,69,66,96,124,81,80,65,
4,3,0,2,5,22,12,23,4,0,0,3,3,67,29,60,85,87,84,84,86,84,83,82,83,80,125,16,81,120,76,76,72,115,93,51,50,76,54,120,149,52,61,73,16,15,44,28,31,34,40,52,71,138,153,114,67,103,151,149,125,159,71,32,32,70,58,87,27,86,119,38,27,32,61,42,29,194,175,182,186,185,132,81,88,93,120,186,186,182,186,189,186,183,221,224,58,11,8,13,13,23,27,26,48,217,214,101,187,183,186,185,185,187,177,186,190,179,187,182,185,187,184,184,184,184,180,185,208,211,13,15,15,15,20,23,21,26,26,221,216,149,180,188,183,186,182,183,186,189,182,187,184,184,187,188,185,192,182,186,184,176,211,217,52,2,11,9,18,45,32,26,93,217,128,177,182,184,187,182,183,179,185,181,175,176,180,177,149,58,79,89,165,196,207,197,194,197,241,221,89,56,67,108,81,62,90,63,59,58,115,122,96,127,122,107,39,42,55,26,122,127,125,123,121,32,11,37,31,46,52,51,83,67,64,63,61,59,135,63,160,102,128,57,136,61,17,88,146,130,185,88,150,69,86,72,
3,1,3,3,14,39,13,11,0,2,9,24,90,86,86,77,85,85,85,82,84,84,81,81,82,79,127,15,76,119,74,75,71,115,84,49,50,49,51,114,71,51,49,36,9,22,28,24,27,18,27,60,56,127,152,105,66,98,97,106,99,82,117,54,68,49,97,70,69,47,67,56,37,23,54,48,50,189,189,191,190,188,67,89,84,100,115,189,188,184,180,191,190,191,231,225,88,96,114,128,145,168,165,175,231,222,219,105,192,186,189,190,186,189,188,185,191,191,188,187,185,190,190,188,189,186,183,191,225,221,54,46,53,47,53,61,52,53,148,219,212,101,183,184,186,190,186,186,190,189,184,189,187,186,190,191,183,194,189,187,180,181,210,213,40,14,15,20,25,26,25,26,75,212,216,101,182,183,184,182,182,180,185,187,183,185,185,182,144,48,79,86,164,223,232,146,193,198,227,231,89,101,78,107,93,53,118,108,38,29,101,118,89,125,124,79,18,46,64,43,124,126,130,129,53,46,36,45,54,66,26,52,63,16,12,119,48,132,132,72,96,95,170,26,80,42,13,94,122,125,157,73,106,99,67,63,
3,2,1,9,8,3,1,6,5,8,7,25,73,83,85,87,86,86,84,83,83,83,83,81,79,79,126,48,68,117,76,74,71,115,79,47,49,50,39,76,50,39,18,14,8,23,14,55,40,44,61,82,64,102,118,144,141,102,123,86,142,98,96,104,55,59,48,53,55,151,26,40,76,36,44,53,154,183,175,176,180,129,180,166,56,79,131,193,190,192,192,196,186,192,219,222,206,218,224,225,220,220,202,222,229,217,219,119,182,185,190,192,193,188,192,191,192,192,189,193,195,196,198,191,192,198,189,189,228,227,201,204,208,185,201,199,194,200,202,162,187,128,185,189,188,190,193,185,193,196,188,196,189,188,193,191,189,189,187,186,183,189,222,219,212,217,227,228,230,224,223,226,227,219,212,106,190,189,188,187,187,189,194,191,193,185,192,186,171,101,76,88,38,170,203,168,192,195,196,209,95,100,101,105,99,34,111,110,103,45,114,102,70,123,122,31,45,49,46,94,102,119,160,126,90,80,88,29,30,24,82,48,91,18,10,111,97,81,75,84,144,80,195,89,98,44,15,112,92,80,94,82,165,128,109,79,
2,1,2,3,2,4,12,13,13,6,22,41,62,35,56,67,86,84,84,83,83,83,83,80,78,70,120,116,118,115,116,73,71,113,74,47,49,47,50,119,28,25,17,9,5,13,14,13,16,53,79,76,82,140,135,148,132,114,124,94,90,70,88,53,58,71,51,78,45,67,49,31,56,56,52,132,139,146,145,142,142,93,102,129,146,151,157,157,155,156,157,156,154,147,148,155,153,155,156,153,164,165,168,166,159,162,162,160,161,164,163,162,162,161,164,157,166,165,169,162,171,171,171,176,186,194,195,196,194,201,197,196,196,195,197,200,198,199,209,210,203,200,203,220,220,221,203,216,214,208,209,215,213,216,215,213,210,197,192,184,176,178,183,182,183,185,177,180,171,169,165,187,197,209,205,126,192,191,192,190,187,192,194,188,181,177,178,189,185,63,67,53,56,40,249,208,192,193,246,216,95,99,102,138,141,131,150,115,52,25,121,99,144,154,125,98,64,51,93,103,62,158,158,160,171,161,139,70,77,40,35,108,32,14,94,50,98,71,74,130,74,83,185,75,78,38,14,94,69,111,65,117,91,151,71,78,
1,2,1,8,9,23,20,29,33,115,28,73,101,81,66,85,85,83,83,82,83,81,82,80,79,70,115,117,116,109,100,73,71,111,54,19,21,21,21,137,16,36,16,7,13,3,13,13,39,46,111,101,104,135,105,156,90,106,122,106,96,61,33,53,47,23,115,132,24,48,75,57,31,27,41,180,136,139,138,137,138,58,106,132,143,144,144,145,148,148,143,146,146,148,146,145,147,143,143,147,147,149,148,152,147,150,148,152,150,149,153,152,149,150,152,153,151,148,152,150,153,142,155,153,153,153,149,151,147,148,147,145,145,143,138,144,143,147,147,148,151,150,152,152,156,160,163,158,148,153,149,150,154,143,161,165,160,156,149,156,147,149,144,135,130,133,143,149,152,153,147,150,143,154,135,136,137,132,136,139,146,146,145,140,140,133,140,137,132,46,94,126,128,132,248,216,158,189,220,225,96,99,102,141,31,33,149,121,97,108,119,85,148,41,61,156,124,72,131,107,53,152,14,55,155,167,143,73,150,106,106,178,86,123,85,45,47,70,65,111,110,110,183,117,53,85,11,73,61,65,70,128,107,130,78,80,
0,27,4,10,18,41,44,21,109,40,77,101,31,109,67,83,82,83,82,82,82,80,80,80,77,71,61,63,61,63,72,72,71,112,49,24,21,24,18,186,12,11,13,9,2,4,12,17,61,26,137,129,162,117,99,119,81,85,83,118,97,71,37,54,26,48,90,94,22,64,141,79,55,21,26,155,157,126,116,134,130,28,90,115,128,127,129,134,135,139,141,141,143,144,144,143,146,150,144,143,151,148,152,150,145,141,147,144,144,150,152,152,152,151,154,155,153,151,153,153,152,146,154,152,151,152,152,154,150,149,147,150,150,152,152,150,148,151,144,149,151,150,150,156,156,153,154,152,151,156,148,149,152,152,151,155,153,158,152,157,143,154,153,150,154,151,149,152,152,148,152,151,152,151,153,146,155,148,148,149,148,143,148,140,137,143,138,131,134,37,71,126,117,127,254,221,132,195,244,225,97,97,144,38,8,10,73,152,115,107,83,154,20,13,9,127,161,39,128,121,146,0,12,19,117,177,144,173,83,133,170,179,166,160,132,141,48,33,74,144,118,130,217,145,65,88,24,19,144,51,87,69,68,68,67,53,
3,132,44,74,22,31,39,58,41,30,23,52,58,35,86,78,82,83,83,82,82,79,80,78,80,74,70,65,70,70,70,71,68,110,44,23,16,18,19,172,14,6,24,2,0,7,14,23,32,47,103,148,136,149,140,92,89,20,64,51,67,75,61,42,13,62,73,59,27,48,135,78,51,73,38,20,64,100,86,69,68,61,38,69,71,74,75,72,76,75,74,74,75,73,75,74,76,81,76,85,94,116,115,84,79,81,82,94,95,114,129,116,103,119,123,135,124,136,131,154,159,156,157,159,156,157,159,158,158,159,160,160,158,158,160,162,161,164,162,163,161,163,165,163,166,165,166,167,167,168,169,170,168,168,168,168,169,168,168,168,167,168,165,163,163,164,165,162,162,161,161,158,156,153,153,153,149,147,142,137,137,140,140,137,138,154,161,153,141,23,129,156,127,83,250,206,190,170,235,189,94,95,129,13,8,6,9,153,115,116,113,152,7,11,4,33,149,39,125,108,149,3,16,9,93,123,129,111,112,84,101,165,192,179,126,180,134,80,132,122,120,98,201,131,80,45,28,18,64,91,66,56,134,104,92,157,
5,106,43,43,48,71,57,42,64,69,78,55,73,51,81,82,84,83,83,83,82,80,79,78,79,74,71,26,59,71,73,72,69,108,35,24,21,21,15,116,15,4,7,4,7,11,14,33,48,69,77,102,142,93,111,80,54,40,46,52,31,71,105,49,78,59,22,47,20,26,122,80,45,57,13,28,52,179,74,75,73,54,27,72,78,79,80,81,81,83,83,83,83,84,83,85,84,84,85,88,86,86,86,88,85,85,88,86,87,86,85,87,89,87,88,87,86,88,88,87,87,88,88,89,89,89,89,88,88,88,87,84,87,89,90,90,87,87,88,89,96,89,88,88,89,89,85,86,87,89,89,88,89,89,87,89,89,90,89,87,87,85,86,85,86,90,87,89,89,89,89,86,86,86,86,87,86,83,84,81,79,79,81,84,82,83,79,100,56,30,67,70,33,48,254,215,216,178,219,211,88,93,126,17,18,16,13,146,116,116,116,149,14,15,16,21,152,53,125,127,153,20,20,29,165,148,100,130,30,40,132,122,118,115,129,124,108,70,91,151,70,80,217,144,107,86,18,17,57,45,82,58,55,127,77,71,
5,72,32,93,68,89,77,76,60,83,81,77,63,86,81,82,84,81,85,83,81,79,78,79,71,63,33,43,31,73,73,71,69,109,39,26,23,16,47,42,13,3,2,7,8,10,14,29,58,43,86,77,97,108,76,95,70,85,89,43,32,55,85,49,47,28,41,63,39,28,123,86,39,33,21,12,32,176,170,81,77,58,33,72,76,80,84,84,85,84,85,85,87,88,88,88,89,88,88,89,87,88,90,88,89,88,88,89,87,89,90,90,90,89,91,91,91,90,91,90,87,92,90,90,91,87,90,89,88,88,90,88,90,90,91,90,89,90,88,89,92,90,89,89,91,92,89,90,92,88,89,90,88,91,89,92,91,90,89,90,89,90,89,88,87,92,92,91,90,91,89,90,89,91,90,91,89,88,89,88,88,86,87,87,89,90,107,144,39,15,78,77,55,40,250,225,130,192,248,223,91,96,99,17,15,15,11,113,113,117,117,115,19,21,20,24,122,58,123,127,124,19,21,35,147,158,115,87,42,47,109,113,112,94,222,77,127,127,72,164,81,101,105,158,112,72,13,17,83,72,100,79,81,112,84,73,
3,16,9,33,71,84,76,73,80,83,82,82,84,83,83,82,83,81,80,82,71,81,79,77,76,42,16,17,38,65,72,72,71,106,41,23,18,11,61,8,11,3,7,3,5,5,10,11,63,64,89,128,75,46,73,70,62,69,57,53,32,50,61,42,60,36,37,44,40,30,134,78,60,32,34,70,83,179,168,168,79,64,25,73,80,82,84,86,86,88,87,87,87,88,90,88,89,87,89,89,88,86,87,89,85,86,89,92,88,91,91,91,91,91,92,91,91,91,92,91,90,91,91,91,92,90,93,92,93,91,93,92,91,92,91,92,92,92,91,92,93,92,92,94,92,93,91,92,93,92,93,93,92,89,92,95,92,95,93,92,92,92,92,93,92,95,96,95,93,94,93,92,93,93,94,93,91,91,91,91,90,90,89,88,92,92,89,84,33,52,78,82,59,40,252,228,225,183,212,223,92,96,99,2,2,2,3,112,112,114,117,116,16,20,12,24,122,71,125,125,123,6,3,26,147,137,152,41,116,89,92,45,83,152,119,151,71,63,127,92,90,94,67,223,137,138,66,17,47,80,88,83,54,169,87,144,
4,7,18,16,72,61,62,53,82,85,84,83,84,86,84,82,85,67,70,42,46,81,82,57,65,15,9,37,58,46,61,65,64,73,44,23,11,9,57,4,2,3,6,5,4,4,28,23,42,81,62,51,125,50,60,50,26,54,28,46,67,68,50,29,35,26,31,61,24,32,88,91,80,31,52,20,51,179,158,174,175,80,27,76,81,84,84,85,83,87,88,87,86,89,91,88,89,88,88,91,89,91,92,89,89,90,92,91,91,90,93,90,92,93,91,91,90,92,94,93,91,92,93,90,90,92,94,93,92,93,93,92,92,93,93,93,94,93,93,93,93,94,92,93,94,93,93,92,91,94,93,94,92,95,94,97,94,95,93,92,92,93,93,93,92,97,97,94,97,94,95,96,93,94,94,93,93,92,92,90,91,90,90,89,92,92,93,86,46,56,82,84,58,43,253,209,158,185,224,211,89,93,97,1,3,4,4,109,111,115,115,115,13,18,10,26,122,68,125,124,123,7,7,62,152,78,135,96,46,28,69,129,80,121,103,66,57,70,85,84,63,72,46,222,132,123,145,16,19,93,102,83,64,89,160,99,
5,10,37,20,20,28,13,48,82,86,84,84,85,80,82,62,49,66,40,23,58,54,67,31,11,21,14,11,69,34,68,78,104,101,49,64,9,8,46,6,1,3,1,5,7,6,8,21,50,55,11,113,126,84,64,91,93,26,46,40,46,35,24,35,28,29,27,31,25,34,165,88,47,139,25,13,7,179,173,171,173,167,37,77,82,82,85,88,88,97,101,108,92,91,117,115,117,109,107,111,117,105,101,103,97,104,110,99,100,102,114,129,129,121,125,110,101,100,102,93,93,93,94,92,92,92,91,95,95,97,92,93,93,95,94,91,94,95,94,93,95,92,95,94,93,95,94,95,94,94,96,105,104,98,96,98,97,97,98,95,91,96,93,93,96,98,97,96,96,96,96,95,94,94,95,94,92,92,92,89,92,92,90,89,93,94,94,89,90,61,81,88,59,43,252,202,124,194,248,215,89,93,97,7,6,4,5,109,110,113,114,115,10,16,9,20,117,73,119,110,101,23,20,87,160,133,98,49,20,159,50,56,79,170,165,135,40,88,68,188,95,144,73,217,130,101,90,24,22,60,121,62,57,45,125,49,
9,10,14,32,56,27,30,63,81,81,81,77,53,78,46,59,64,36,12,16,19,45,14,12,8,5,4,24,44,145,101,88,42,55,37,22,7,14,6,4,4,7,0,37,1,4,10,6,8,12,38,84,131,71,61,84,60,39,22,30,58,24,18,34,23,21,27,27,15,30,176,85,36,144,31,20,10,168,170,173,173,175,29,77,84,85,86,180,93,89,179,184,167,91,91,173,172,178,177,176,177,181,175,182,178,179,183,178,178,181,185,182,179,179,172,182,173,191,170,183,179,174,183,184,180,181,183,180,178,183,178,179,175,179,186,180,185,181,179,175,183,180,177,179,182,182,179,183,179,183,192,181,177,180,177,182,183,182,187,187,179,184,173,183,180,181,183,178,181,175,163,179,183,161,150,142,124,99,96,96,97,92,90,94,102,116,162,181,148,62,85,88,42,53,253,203,213,189,222,217,82,91,95,2,5,2,6,106,109,111,113,115,10,21,10,16,118,83,120,122,121,7,7,145,146,160,60,29,6,14,113,122,47,98,134,80,82,47,125,74,93,74,177,205,99,82,145,40,21,51,61,42,194,124,64,66,
9,9,15,12,16,8,18,72,70,77,65,43,36,58,16,59,22,17,8,13,12,11,8,39,61,4,17,39,57,40,33,57,62,56,42,14,9,6,6,5,4,3,3,3,3,11,6,2,16,37,58,57,110,73,84,22,58,15,31,16,49,22,21,38,19,36,36,23,15,24,172,77,26,39,19,19,16,170,175,173,168,182,26,77,82,85,88,176,176,154,90,120,167,92,93,100,174,174,176,179,175,179,173,177,176,177,181,178,181,181,189,181,178,176,174,179,178,177,172,184,181,177,184,181,182,178,179,180,179,178,176,181,174,180,180,181,181,182,180,181,179,181,178,182,181,181,179,183,182,180,187,182,182,183,180,187,186,181,184,177,168,180,181,175,174,180,181,185,183,187,179,183,185,180,184,184,178,177,182,175,183,174,175,178,179,188,184,181,148,62,86,88,6,17,253,218,150,193,245,228,82,88,93,1,4,1,5,106,105,107,110,112,12,21,10,17,115,80,115,118,120,4,7,85,174,113,78,105,29,27,61,75,72,94,120,47,67,50,41,74,53,60,136,122,105,84,161,42,22,32,28,43,168,51,140,82,
7,4,4,16,6,12,34,74,96,99,70,43,75,41,47,10,33,11,4,6,8,6,5,8,13,2,3,12,44,30,29,43,36,89,51,9,11,1,1,1,2,2,5,4,3,20,46,53,50,95,122,68,92,92,66,26,45,45,16,37,54,44,18,24,12,45,46,20,15,25,197,69,25,59,17,12,15,177,180,173,176,179,27,78,83,85,90,177,178,176,175,92,87,89,92,90,162,175,173,177,178,178,178,179,178,181,184,180,180,182,185,180,176,175,181,180,179,181,178,180,178,178,188,179,176,174,177,178,180,178,179,179,180,177,182,181,177,179,184,182,180,180,174,181,180,182,181,173,180,184,183,180,184,181,184,182,182,185,183,175,177,179,172,179,181,183,185,186,181,183,178,183,182,179,186,181,179,178,180,179,179,177,178,180,184,182,183,186,143,63,85,88,21,17,253,185,169,191,227,199,80,85,91,7,8,6,7,102,103,104,107,110,9,17,16,18,110,86,109,111,117,12,6,20,156,133,143,28,70,45,28,51,95,62,128,95,111,72,37,81,53,182,82,82,190,140,123,41,23,20,45,70,157,66,62,85,
5,5,5,10,9,44,88,138,135,106,53,62,37,42,45,8,14,5,3,9,4,2,13,7,3,3,3,7,25,13,37,41,18,70,17,7,5,2,1,2,9,5,9,10,6,34,44,43,31,59,75,44,60,119,69,40,24,27,18,43,82,39,20,8,5,45,44,20,13,22,154,62,29,54,13,13,26,177,177,173,176,179,30,77,83,85,88,179,178,181,180,182,96,88,88,88,90,175,178,176,177,174,182,178,177,179,182,176,178,172,183,182,174,181,174,174,180,187,183,184,177,178,183,181,177,179,180,178,180,178,178,181,177,180,181,180,174,185,181,187,177,179,180,180,179,179,184,173,181,177,183,180,183,184,184,175,186,185,180,173,173,180,177,181,178,183,184,184,179,176,176,183,185,184,188,184,181,176,176,182,178,179,177,180,178,175,184,184,141,53,86,89,112,125,186,209,227,200,218,215,96,107,108,105,105,103,110,117,118,121,120,126,114,115,112,116,133,92,124,83,126,22,25,44,176,128,54,62,69,31,89,49,158,126,140,104,106,74,71,54,60,96,112,105,210,129,164,52,64,63,56,59,77,23,140,159,
10,4,8,14,15,105,117,136,132,118,56,26,33,21,10,10,7,3,8,4,8,2,1,66,2,2,4,13,72,33,20,40,10,29,18,15,35,3,1,3,4,5,24,15,10,14,37,77,44,71,29,23,51,46,28,44,33,15,19,36,34,25,15,17,5,48,44,18,10,21,162,25,37,56,16,13,49,179,178,177,175,180,29,78,85,85,87,178,174,176,179,180,181,146,89,89,91,168,175,177,178,179,177,176,180,171,178,176,180,174,181,180,173,179,174,175,179,183,181,172,181,180,183,179,180,179,179,180,182,181,177,179,181,179,179,172,176,176,181,174,177,179,181,178,181,181,184,184,187,182,177,181,180,184,178,179,183,187,183,174,177,179,179,185,177,178,185,180,179,178,179,179,180,180,183,184,176,174,177,180,177,178,177,183,178,179,181,182,138,63,86,88,165,181,136,156,206,206,208,210,33,31,33,34,36,37,38,41,40,43,43,45,44,49,81,127,151,92,124,104,116,23,28,71,159,138,76,17,21,17,121,41,78,107,64,79,35,61,45,80,89,66,77,104,202,93,151,69,55,21,58,124,117,112,81,89,
8,3,13,15,68,110,102,111,117,125,70,60,15,9,16,12,7,7,8,4,2,3,8,2,10,8,6,7,115,38,24,34,12,22,39,56,58,3,1,3,53,7,0,4,18,65,152,154,74,43,27,68,42,18,33,14,13,17,16,22,27,28,25,23,8,49,41,16,11,18,182,20,57,57,11,36,72,167,174,176,179,177,29,79,83,86,88,177,172,177,182,180,183,182,174,151,117,166,170,177,178,170,178,179,179,180,179,180,180,180,186,182,171,180,172,185,185,179,178,175,176,178,185,180,178,178,180,178,180,178,171,174,180,186,214,165,176,176,183,174,181,184,183,179,178,183,184,183,184,179,186,181,182,183,181,178,178,184,182,168,176,176,182,182,175,181,183,177,175,181,180,179,176,178,185,183,180,183,178,185,181,180,178,180,179,176,184,183,140,64,87,90,86,118,89,76,69,86,73,84,32,31,31,34,37,36,39,42,38,41,41,45,45,108,63,160,143,95,120,35,40,137,26,84,171,150,117,68,57,13,80,74,20,13,16,111,93,68,51,56,62,46,129,135,196,98,172,81,39,28,119,93,142,75,59,70,
6,3,8,11,67,130,107,75,77,73,45,23,14,11,1,2,1,6,5,4,3,1,4,14,1,6,5,69,223,32,17,24,16,21,35,31,4,23,12,3,11,40,64,113,158,91,108,184,101,124,37,65,67,47,46,26,53,20,16,18,20,19,24,21,9,66,46,16,64,41,172,48,29,66,15,58,17,180,174,176,183,173,27,79,83,87,89,178,173,181,186,179,173,178,173,178,168,179,171,231,165,93,176,181,175,180,175,178,177,182,178,178,173,181,178,184,177,183,179,175,179,180,185,179,176,179,177,177,180,174,173,173,179,216,238,118,152,181,183,179,176,182,182,178,178,185,184,186,178,178,184,179,180,177,183,179,183,190,183,172,179,181,181,180,173,180,179,243,214,221,176,177,177,181,187,180,182,181,178,188,179,179,175,181,180,179,186,182,132,63,88,89,135,132,93,133,74,75,84,144,29,27,30,33,34,35,36,38,34,37,40,40,41,216,217,204,216,105,33,24,30,18,11,135,164,72,57,103,76,17,28,26,9,14,91,53,48,22,57,74,45,61,61,43,118,91,157,89,77,33,29,52,56,112,69,102,
5,3,11,18,19,65,80,77,79,78,15,20,2,1,0,2,1,1,3,4,2,3,7,18,23,12,105,78,127,61,11,17,34,53,33,7,13,64,10,3,48,28,167,107,89,83,133,120,108,69,51,62,70,42,32,18,60,40,49,14,13,52,67,72,155,186,173,77,77,84,183,28,124,177,64,68,12,153,178,181,186,177,29,78,83,87,88,176,172,172,177,178,176,174,173,179,169,178,180,243,155,83,92,174,178,174,175,175,172,179,181,180,180,181,180,183,182,175,179,178,181,185,178,181,181,179,176,178,176,174,172,176,178,236,211,116,78,156,176,178,176,182,181,182,176,182,181,185,177,182,181,181,181,180,181,175,178,187,180,170,175,182,180,182,173,175,176,239,186,152,94,180,182,181,180,185,181,180,178,184,179,179,177,180,184,181,181,184,130,63,87,89,65,129,104,127,144,98,69,113,35,36,43,41,47,40,46,46,52,49,53,58,55,212,220,228,226,100,150,89,81,99,60,115,153,157,148,78,23,12,50,48,5,2,63,93,155,92,103,60,121,37,19,90,92,167,116,111,91,36,19,120,82,115,67,116,
4,4,7,5,22,73,77,76,77,76,16,5,16,4,4,1,4,2,2,1,5,9,10,50,17,53,101,57,58,57,20,27,26,51,1,29,17,23,20,16,8,55,79,64,123,132,126,98,113,99,42,122,65,38,33,21,59,70,18,17,19,21,47,116,178,143,135,163,163,186,172,29,167,185,166,162,36,94,117,177,181,179,28,78,83,86,89,174,178,177,177,176,173,174,176,177,190,214,217,249,152,137,143,145,187,171,176,176,175,181,183,184,176,179,177,179,177,178,182,178,179,182,179,172,176,172,177,183,175,175,205,220,214,237,125,121,124,115,93,178,181,186,184,185,182,184,180,187,176,180,183,178,181,181,179,174,175,186,177,172,176,178,184,181,178,174,180,240,169,153,89,96,175,177,181,184,176,177,178,182,185,179,173,181,183,179,179,183,128,61,86,88,168,169,172,191,186,189,189,195,200,198,199,200,197,194,195,194,194,194,198,199,204,226,138,210,241,96,156,158,152,71,210,193,172,155,79,55,45,30,163,79,2,7,38,123,90,99,76,31,69,37,47,112,104,72,132,119,121,87,22,65,128,75,149,52,
3,10,3,17,25,8,5,7,3,8,4,9,4,3,1,2,1,0,1,6,8,2,6,49,20,58,88,4,17,13,5,14,13,3,7,22,43,11,8,44,90,36,33,73,58,89,101,80,39,53,73,58,28,41,47,13,27,28,99,63,22,15,67,98,122,115,75,121,146,191,197,25,139,133,136,179,76,86,90,130,175,176,28,80,84,86,91,175,177,186,176,175,179,178,183,221,213,222,221,246,144,144,150,223,220,215,214,151,175,179,183,183,176,179,172,178,181,183,181,176,177,176,178,177,177,171,179,180,174,222,215,222,217,225,151,129,136,137,138,176,177,181,184,186,182,184,179,189,178,182,181,178,184,176,184,179,174,183,178,173,172,182,180,181,187,222,222,245,162,148,150,222,181,176,177,183,178,176,182,180,185,178,178,180,179,180,178,181,128,63,88,88,207,213,209,210,211,210,210,208,207,204,210,209,207,206,205,212,206,209,207,206,206,152,214,214,149,103,174,156,135,135,204,206,166,162,39,22,59,34,96,16,4,23,53,50,127,99,90,69,100,49,48,135,12,166,146,153,136,104,28,26,48,80,65,102,
1,2,2,1,7,28,54,75,93,1,4,13,22,9,1,4,4,1,23,8,4,21,47,159,60,58,63,5,16,41,11,14,4,7,30,24,16,18,12,49,70,33,31,67,107,97,85,61,66,52,56,84,34,28,76,61,63,145,121,92,53,14,27,54,37,44,28,49,57,65,119,38,37,72,86,80,47,91,90,101,146,172,27,79,85,86,93,178,175,183,170,179,187,213,195,153,217,216,150,113,53,33,97,226,210,246,160,89,164,173,178,181,177,179,179,176,179,185,178,178,181,175,181,178,176,181,181,196,218,214,220,210,210,169,58,97,120,126,130,139,228,210,174,181,183,182,179,184,176,178,184,175,186,211,210,212,207,178,175,173,175,185,182,212,215,219,222,222,157,154,150,222,221,214,194,179,178,179,179,180,183,182,180,182,179,173,178,182,125,67,88,88,206,206,206,207,208,207,209,207,207,204,210,185,168,175,185,191,179,171,173,173,178,125,49,41,181,105,127,110,125,101,75,152,158,82,96,35,29,11,122,4,6,58,29,29,161,46,45,55,17,44,119,5,11,166,82,158,165,147,96,42,40,35,100,90,
2,1,1,7,25,59,75,115,130,121,70,31,12,44,7,4,3,3,4,23,34,46,34,107,61,61,61,4,8,33,12,3,5,17,19,34,28,64,55,34,84,31,63,91,77,64,116,37,21,25,53,53,25,37,50,36,78,68,116,70,31,19,28,26,20,44,22,31,40,92,62,16,99,40,62,31,30,89,89,86,107,135,22,79,85,87,98,182,185,179,173,178,181,220,164,145,40,21,23,16,19,25,24,27,29,168,161,86,86,177,178,179,174,179,175,178,177,183,172,175,179,170,179,176,169,182,183,224,161,211,126,34,25,7,18,30,8,12,39,116,141,140,94,182,182,177,173,185,181,176,178,174,223,25,21,24,29,220,172,173,176,193,231,167,216,143,27,24,22,21,29,108,224,248,165,85,181,177,179,175,181,177,176,179,179,179,177,181,118,65,89,89,205,204,205,205,207,207,208,205,207,205,205,205,206,208,189,197,207,194,208,200,182,194,188,201,110,112,15,15,23,10,30,36,136,169,102,29,9,8,26,5,5,109,34,22,188,10,88,154,98,65,82,4,14,153,114,177,131,162,49,18,60,37,109,9,
1,5,0,10,16,22,49,131,129,124,44,10,44,32,3,17,5,22,10,16,8,36,52,93,64,50,19,5,6,4,9,2,10,18,24,27,16,36,18,44,49,36,36,77,80,82,46,35,21,36,38,38,36,39,63,67,114,84,96,51,40,25,22,18,17,18,23,28,37,45,26,17,62,53,37,26,9,101,84,86,97,84,23,79,85,86,101,181,178,172,173,182,183,226,156,157,20,5,7,25,45,49,31,20,30,176,164,83,88,165,178,180,175,181,178,174,178,185,181,181,181,178,178,174,177,176,186,230,176,33,9,18,29,6,49,28,25,7,9,34,127,155,89,122,182,178,173,187,186,177,177,174,227,14,10,8,10,212,96,173,177,194,188,169,28,27,26,19,40,20,15,27,34,190,140,81,94,173,179,177,181,180,178,180,177,178,178,179,115,65,89,89,204,209,206,208,208,209,203,206,210,206,205,205,204,205,209,205,210,192,219,201,206,212,204,198,206,86,204,208,197,197,195,203,175,162,89,23,19,21,27,1,25,106,10,73,160,23,126,103,66,60,99,42,3,125,146,160,164,114,42,27,29,61,24,48,
6,8,0,9,6,45,36,132,11,6,54,24,28,21,38,24,8,12,20,51,39,32,33,47,63,60,44,3,5,7,0,17,26,28,39,26,27,25,25,24,37,44,46,19,60,72,28,11,30,30,46,45,42,39,50,42,61,71,56,31,60,27,21,11,21,17,22,34,18,29,59,6,49,41,19,21,5,90,124,84,94,81,23,79,85,87,104,179,176,177,172,179,178,226,158,148,19,2,8,27,26,66,99,34,25,203,148,83,91,165,181,181,170,179,174,177,175,176,176,179,181,175,172,175,177,182,186,219,163,34,13,7,25,7,19,31,53,11,7,33,79,152,91,119,137,120,138,138,179,180,181,171,218,12,11,6,11,215,94,174,178,202,161,166,18,14,15,68,58,11,33,16,32,177,158,83,96,178,178,180,182,181,181,180,176,175,180,180,116,66,88,89,206,205,205,205,206,203,205,203,203,204,205,202,201,198,198,197,197,200,189,196,205,221,217,195,198,111,217,214,205,214,216,217,156,129,134,24,12,13,2,5,31,96,9,44,206,14,83,118,51,59,93,66,10,14,161,164,172,98,120,26,36,46,46,79,
37,16,12,8,7,66,76,131,19,9,50,53,50,35,49,42,17,53,38,36,49,60,65,59,63,61,31,2,2,2,26,11,5,13,10,15,28,33,47,17,26,24,31,51,20,17,6,18,37,74,27,44,31,35,35,43,46,59,68,35,22,37,31,44,22,30,24,19,43,81,44,8,71,10,12,17,1,89,85,86,85,73,22,78,84,86,98,161,177,184,173,180,176,179,118,143,16,3,6,21,28,35,49,98,25,196,199,86,89,167,179,178,167,183,178,174,177,176,177,178,178,178,180,177,179,184,178,209,144,33,20,8,27,11,16,32,12,10,9,36,153,158,87,125,135,98,141,141,114,180,176,173,217,12,8,12,13,213,92,174,179,197,160,164,17,7,9,35,49,72,33,15,31,192,156,87,94,178,178,178,180,181,181,181,178,179,182,180,111,66,88,90,206,202,198,202,200,197,201,199,198,198,200,199,197,201,202,202,204,201,202,200,193,200,198,207,209,120,209,204,207,211,215,205,166,126,120,41,52,87,62,17,75,21,44,18,164,35,110,101,78,65,33,61,11,59,155,183,171,114,24,29,45,32,65,36,
16,9,5,9,8,63,78,130,18,10,28,37,97,58,38,41,34,14,45,52,50,61,62,62,63,59,55,0,1,13,27,15,3,15,7,73,12,37,22,16,34,14,16,24,18,6,6,15,48,43,28,42,35,22,48,59,40,35,34,19,27,18,31,25,31,16,23,34,42,68,4,28,50,20,19,40,7,87,101,84,93,65,21,79,84,86,89,127,146,174,167,180,177,171,230,217,14,25,16,11,16,19,22,54,20,210,194,123,162,174,181,177,168,179,177,175,178,177,181,184,183,181,175,174,181,184,169,232,184,33,19,14,28,10,14,33,10,5,7,36,140,150,87,139,128,77,130,134,132,146,176,177,218,6,3,2,10,215,93,175,180,181,135,154,16,8,41,79,74,78,44,13,39,224,122,94,95,178,175,180,180,184,176,181,178,176,179,182,111,65,88,90,203,199,201,204,210,217,219,215,209,198,195,194,194,193,194,194,193,195,198,200,203,202,208,203,210,162,182,179,181,184,188,194,166,145,124,114,122,117,149,102,141,121,28,21,193,53,36,48,120,129,137,63,17,72,187,168,182,143,82,31,19,72,22,33,
66,37,25,4,6,43,76,130,14,6,32,27,69,57,45,60,58,52,50,65,27,31,17,26,5,5,3,1,2,50,34,5,4,8,8,38,19,12,8,34,34,7,21,19,27,3,16,15,21,84,41,34,50,30,46,48,48,20,21,13,43,17,27,23,24,29,23,35,50,14,37,28,31,10,3,6,102,111,93,91,82,71,21,79,84,86,88,110,104,104,156,181,180,171,223,211,14,17,16,21,22,23,60,39,22,215,188,148,174,164,178,179,173,179,186,178,176,175,181,182,177,174,175,176,176,181,171,232,205,44,24,18,28,11,15,31,8,10,11,37,140,153,95,128,121,96,109,131,92,169,179,175,223,5,1,0,5,214,94,175,178,176,217,214,32,23,25,23,38,25,26,29,49,223,149,94,97,180,175,177,181,181,176,179,176,177,180,180,111,65,88,90,176,209,207,204,206,208,210,210,210,204,191,203,193,193,195,193,192,190,192,190,193,200,198,200,200,200,201,199,197,198,156,172,168,141,99,107,107,88,164,88,84,88,76,187,189,185,98,75,124,175,70,193,9,32,199,149,181,124,130,85,21,51,48,192,
75,29,21,4,2,12,76,128,16,9,35,55,110,47,68,69,70,67,65,24,9,2,4,4,4,24,49,3,8,2,2,7,2,14,16,6,16,8,60,14,5,6,18,9,2,3,4,33,24,33,26,26,21,25,59,103,45,36,16,23,67,36,16,23,18,23,32,62,37,15,11,6,18,9,6,62,9,123,108,95,88,68,21,79,84,86,87,116,102,95,95,147,178,159,219,213,43,41,45,50,55,17,12,15,66,212,188,155,171,164,174,182,171,182,176,177,174,180,182,178,174,175,175,174,176,176,170,231,205,43,73,75,47,72,14,55,63,80,97,37,143,154,95,182,92,97,101,98,99,176,180,177,219,4,1,1,8,214,96,172,177,174,215,215,16,8,12,33,59,32,18,15,27,215,149,177,179,179,175,183,181,182,180,178,178,175,181,181,109,67,87,89,210,210,209,208,208,206,211,210,208,206,204,204,198,220,205,192,204,202,202,206,199,199,203,199,207,200,207,209,203,194,168,110,125,147,130,159,151,65,95,105,57,100,68,107,80,132,90,32,42,176,53,35,14,14,213,142,203,151,182,86,26,103,48,37,
13,12,11,3,2,12,57,89,11,6,40,61,121,66,67,65,63,14,2,1,3,6,18,21,52,59,50,2,13,15,3,3,1,10,1,4,4,4,6,1,10,10,4,1,2,1,3,14,14,68,24,38,32,36,30,41,46,42,26,39,107,50,30,59,46,17,42,4,19,8,5,5,65,15,3,155,5,101,118,111,83,68,19,79,85,86,99,117,104,99,106,92,144,171,210,193,17,4,7,11,20,42,52,33,23,200,190,137,179,175,174,184,169,177,178,174,179,183,176,179,177,179,176,173,175,174,172,234,202,40,74,80,50,83,15,58,70,92,108,38,141,151,96,186,142,138,138,129,152,181,174,172,217,5,1,4,8,216,93,171,178,177,212,215,14,8,12,15,18,9,10,10,37,217,158,181,177,177,176,182,181,179,174,171,177,174,177,179,105,65,88,89,158,208,204,208,208,205,202,204,207,207,207,206,206,209,201,199,213,204,206,211,203,204,208,200,206,202,203,211,201,207,208,208,211,173,123,138,161,134,140,162,134,171,151,141,144,157,146,148,139,150,101,83,137,95,156,148,173,173,149,62,27,29,66,33,
14,10,3,3,1,6,15,125,8,4,42,66,120,68,64,3,2,1,1,29,25,8,5,36,52,55,48,4,17,61,7,3,1,1,2,4,2,6,1,3,33,9,2,1,3,2,3,3,6,16,38,34,38,29,46,22,43,35,29,34,110,19,70,97,36,86,28,26,16,8,9,23,36,14,10,113,5,86,127,99,93,71,18,79,83,85,88,141,121,101,110,94,93,131,214,170,16,4,8,10,22,48,53,50,20,210,187,135,174,173,177,181,172,181,174,173,179,182,178,179,182,182,172,173,176,180,179,236,205,42,72,76,46,79,15,56,77,97,109,40,144,154,95,130,109,123,127,137,135,183,173,178,217,3,0,2,8,213,94,176,183,172,213,216,17,11,23,26,45,72,48,11,36,220,150,168,181,178,175,183,182,176,172,179,174,173,176,178,105,67,86,80,186,130,205,200,206,205,207,206,208,206,199,199,203,201,202,201,203,201,200,221,211,196,203,198,204,196,183,186,184,190,193,192,194,205,203,208,184,78,158,126,197,145,127,142,144,150,156,173,138,170,198,171,155,142,120,167,192,184,173,99,24,17,77,17,
10,16,16,4,9,4,13,77,17,5,48,65,58,4,2,0,6,16,16,1,1,2,32,42,46,53,12,4,21,20,6,0,2,1,3,2,4,4,3,1,2,1,27,10,9,12,38,19,46,27,9,24,48,56,40,27,24,38,17,63,131,36,12,8,14,22,2,24,52,6,0,4,6,23,14,99,3,85,95,116,97,87,20,78,84,85,89,116,148,126,97,98,88,87,167,182,17,1,9,23,21,49,48,53,22,204,184,121,165,172,175,179,179,176,177,172,181,179,181,178,176,174,170,168,175,180,181,227,206,41,28,26,27,33,19,36,32,44,49,41,158,154,94,122,108,138,132,139,136,115,180,174,223,3,1,2,10,212,95,170,173,170,221,211,20,20,62,27,44,62,59,63,33,228,143,170,174,179,183,183,180,177,175,179,178,169,181,177,104,67,87,124,105,101,86,133,146,153,180,182,173,138,158,146,154,172,185,177,174,190,195,199,195,199,197,172,191,201,192,181,181,205,209,208,207,208,209,214,216,221,212,195,156,149,151,92,147,90,150,188,153,166,129,165,155,176,147,165,142,96,188,148,97,18,158,143,
13,41,5,4,27,2,4,72,18,2,43,5,3,1,22,11,8,1,4,0,3,6,19,20,29,21,12,5,20,58,4,7,0,1,1,2,2,1,0,1,4,4,20,6,10,7,25,37,62,55,49,36,19,24,23,24,20,23,17,27,169,17,77,40,12,7,11,23,9,4,22,6,8,12,18,79,4,84,87,96,95,99,21,77,85,86,87,117,144,149,110,92,87,85,122,160,16,32,54,50,22,45,43,55,22,211,183,103,169,172,175,178,175,177,177,177,178,180,178,175,174,167,171,173,173,173,171,226,78,27,16,16,24,17,16,30,18,17,19,40,172,152,93,135,140,138,140,137,94,173,177,174,228,20,21,23,33,218,93,175,178,172,221,216,30,18,50,28,43,70,59,57,32,223,149,164,173,181,183,177,178,178,176,177,179,175,178,177,98,67,88,73,209,227,36,61,66,61,60,55,55,54,55,57,57,56,56,59,57,57,57,63,90,79,87,92,191,175,195,188,176,133,178,170,185,184,173,186,206,208,209,212,216,211,203,168,155,96,72,97,62,102,163,184,139,155,144,108,22,26,34,60,74,21,54,98,
42,76,7,9,23,2,6,84,15,6,1,2,54,48,41,51,11,4,1,0,8,8,13,15,12,23,10,8,7,51,2,8,2,1,2,3,3,1,3,2,9,18,49,27,6,18,20,22,18,17,11,13,14,18,31,23,17,5,4,6,182,11,9,7,18,16,6,12,62,9,11,6,33,34,3,60,6,83,83,86,85,78,18,77,85,87,86,88,118,137,125,104,91,84,131,148,16,33,54,47,19,47,38,55,21,211,183,103,174,176,184,176,170,173,180,174,182,173,179,173,103,100,87,92,84,75,73,106,81,57,19,14,19,20,19,18,21,22,26,17,151,151,94,183,117,119,119,110,118,178,183,180,228,114,131,149,160,223,93,173,175,169,224,200,36,19,51,26,44,68,57,55,31,218,132,143,180,180,179,173,178,177,174,177,180,175,179,176,99,67,88,78,187,225,37,66,75,65,65,53,54,56,58,61,77,91,94,106,91,83,91,82,79,71,61,74,85,59,89,45,74,55,63,70,59,55,76,72,58,68,80,75,74,72,63,82,73,55,28,76,57,137,93,142,151,105,98,93,18,13,18,24,31,24,43,118,
15,27,14,8,10,2,2,27,13,2,2,37,69,52,27,37,6,5,4,3,5,6,9,29,17,17,6,3,3,8,7,6,4,2,1,2,4,7,4,6,7,66,61,24,12,26,18,31,4,6,16,14,13,12,17,38,103,84,147,103,120,42,8,38,97,111,106,77,75,15,8,12,104,5,9,65,4,83,84,83,81,68,16,78,82,85,87,87,88,108,114,105,95,91,150,151,12,24,48,47,16,44,34,53,20,223,185,105,173,176,183,173,173,175,181,180,179,171,173,171,172,172,89,167,175,162,138,230,202,42,26,21,21,23,25,23,22,29,33,31,146,153,93,165,137,106,102,139,150,182,181,180,235,202,210,218,216,205,95,170,171,168,229,193,31,16,48,25,49,72,59,56,31,224,136,174,177,177,178,173,175,173,178,180,176,172,181,177,100,69,89,76,215,208,55,43,52,52,57,64,68,64,72,69,54,61,64,58,68,70,55,64,55,56,60,68,63,60,55,59,61,52,51,63,61,63,66,59,64,105,136,183,199,202,199,206,204,203,208,208,203,159,90,173,146,144,127,48,16,18,23,27,27,22,20,97,
1,7,3,7,8,6,2,2,1,4,18,22,42,53,12,45,13,11,0,3,2,3,3,13,7,3,6,1,0,8,4,4,5,2,2,4,2,9,17,32,15,19,52,24,24,38,24,24,96,9,2,10,9,7,8,84,90,32,82,98,28,62,3,91,92,73,70,139,65,104,102,156,125,67,69,98,7,85,84,83,82,67,16,77,82,85,90,89,87,90,103,102,107,89,158,166,25,29,36,53,55,29,23,33,117,218,185,111,173,175,174,178,173,179,180,179,178,177,178,175,172,170,87,166,182,172,138,214,204,47,32,21,23,26,29,23,24,31,39,52,144,156,96,139,139,100,84,141,134,182,180,184,224,175,191,210,208,218,97,121,174,176,230,200,37,16,44,24,48,79,58,58,31,218,127,176,176,176,176,163,180,182,181,179,178,176,179,179,99,68,89,71,216,229,182,80,66,117,81,97,108,78,64,78,62,52,55,54,51,54,54,56,57,55,52,52,48,50,55,53,61,59,61,69,55,163,196,204,198,201,201,202,205,209,204,209,208,209,210,208,208,217,215,210,185,187,74,40,21,17,16,28,27,24,20,159,
113,24,11,5,2,2,2,1,2,19,20,19,28,46,4,14,9,2,6,1,2,3,6,15,5,8,5,1,3,0,5,3,1,24,35,7,2,18,9,16,30,33,35,10,23,15,22,10,25,7,1,7,8,6,13,105,60,20,38,39,5,1,10,20,57,35,38,59,47,15,125,115,106,117,63,129,14,85,85,84,82,67,17,77,83,86,86,87,88,91,87,97,100,98,136,153,16,17,15,15,15,45,36,51,22,215,188,113,180,175,173,179,177,177,184,179,181,186,179,173,168,169,94,78,79,75,77,109,119,35,30,19,22,28,29,24,30,32,45,58,140,157,92,141,135,146,143,146,125,97,180,178,167,147,105,101,99,99,98,127,179,180,228,207,24,27,28,23,16,21,27,26,34,217,131,171,175,173,180,179,181,183,182,179,180,174,179,181,98,69,88,69,227,196,126,43,45,209,207,205,210,207,202,202,196,194,195,195,198,195,190,195,201,199,199,202,200,193,200,201,203,200,198,208,194,197,190,209,170,172,206,191,175,202,198,203,209,200,207,207,207,214,205,208,205,208,199,165,21,19,18,25,18,17,22,40,
63,76,22,16,7,3,1,0,1,1,12,14,30,10,8,7,8,4,1,19,5,9,3,6,0,4,0,1,2,2,7,4,5,5,10,6,5,4,8,32,20,90,56,5,3,9,6,6,31,3,6,3,12,6,20,67,35,7,17,114,19,2,6,40,14,54,36,70,52,19,66,83,106,84,117,154,16,85,86,85,81,68,16,77,84,87,86,88,86,88,88,87,101,97,155,151,14,28,49,50,14,46,29,51,17,211,189,104,177,181,175,177,182,180,173,177,183,167,176,172,169,171,91,76,79,73,68,112,121,35,31,22,23,29,30,26,30,35,49,59,137,158,100,146,144,130,123,142,95,174,186,175,173,182,178,182,182,184,184,178,176,180,233,208,44,16,52,29,53,72,55,61,42,219,128,152,176,176,181,183,182,173,183,179,179,179,179,178,98,69,88,77,217,224,156,174,125,203,201,206,200,204,204,207,205,204,204,202,199,201,201,195,193,181,163,134,114,123,105,99,150,173,189,197,197,206,199,194,192,198,217,212,203,207,200,200,200,205,207,213,206,211,211,209,207,203,199,88,21,19,16,15,20,24,19,30,
104,56,40,9,0,10,4,3,9,7,14,20,35,3,9,3,7,8,18,5,8,31,4,2,2,1,1,1,1,1,1,2,2,9,11,8,46,9,4,11,16,30,19,8,5,9,5,4,7,5,3,9,24,6,12,9,8,6,23,18,2,1,6,6,28,20,62,49,31,58,17,52,23,69,25,196,22,91,88,86,81,70,18,76,83,86,85,84,89,86,86,85,103,105,152,154,15,27,53,50,15,46,32,49,18,202,187,98,177,173,172,177,176,181,172,174,186,158,174,176,165,174,90,76,82,71,65,159,114,35,34,22,24,30,32,25,29,37,54,59,141,157,97,185,149,155,156,121,108,182,179,179,182,185,178,184,181,179,179,180,171,173,236,208,41,15,47,30,51,77,54,56,36,221,124,168,176,167,181,181,185,172,184,177,174,176,182,178,95,70,90,74,208,213,205,56,199,201,202,198,202,200,202,201,200,200,202,202,202,200,201,202,201,199,197,196,200,200,196,199,195,196,193,193,197,193,192,198,196,193,190,189,195,216,206,201,201,194,195,202,199,205,206,203,208,204,201,23,25,12,8,19,27,23,17,20,
99,71,35,6,1,2,2,3,2,12,17,7,4,7,6,7,9,25,20,9,35,25,8,7,3,3,1,1,1,2,2,2,4,8,7,5,4,6,9,4,16,20,6,6,7,5,5,3,7,7,8,8,10,3,11,22,12,11,47,6,2,3,3,3,5,33,81,109,44,58,10,39,14,110,117,183,16,85,91,83,83,68,16,77,82,84,84,84,85,85,85,85,88,104,178,146,14,22,50,52,15,47,31,51,17,169,170,102,177,176,177,170,176,176,169,179,182,175,178,173,135,132,86,88,86,82,87,119,103,35,35,21,25,28,32,24,30,37,57,62,140,156,99,112,107,106,103,99,116,180,179,180,181,184,182,180,178,176,177,174,172,174,238,208,42,12,49,29,53,83,60,57,37,222,138,169,174,179,180,180,184,179,177,177,175,181,180,175,93,71,90,74,233,225,170,122,192,177,200,201,199,202,202,199,198,197,199,198,200,202,202,200,200,201,199,198,196,195,198,202,192,196,193,195,193,191,193,192,192,197,202,197,189,187,191,209,217,202,196,196,198,204,198,169,180,172,189,13,17,22,16,18,17,20,13,12,
127,62,12,6,1,2,2,2,4,7,14,3,6,2,4,9,5,19,17,25,13,21,16,3,15,13,7,3,8,4,0,8,3,4,29,17,5,10,7,8,8,28,7,5,14,2,8,3,3,3,41,7,7,6,6,5,3,1,2,5,3,3,2,8,27,21,28,26,13,26,9,16,14,89,42,85,39,84,86,87,82,70,20,77,82,84,84,84,85,85,84,85,87,83,176,174,16,22,55,57,14,46,32,51,14,149,153,114,176,176,183,172,178,177,174,181,177,173,179,176,173,179,99,73,74,70,75,162,123,32,34,23,25,28,32,28,30,37,67,62,139,155,93,104,91,82,97,106,94,182,175,181,181,186,182,181,183,179,180,169,171,174,241,209,46,18,46,28,50,80,58,59,38,220,143,124,179,180,181,184,183,176,178,175,178,181,177,174,93,70,89,73,113,223,45,49,62,49,56,66,52,90,196,200,193,198,197,197,199,200,199,200,203,200,202,202,200,198,199,196,196,199,197,199,198,196,196,193,192,190,193,197,197,194,197,191,185,176,87,40,47,47,43,47,61,80,18,20,19,21,13,16,14,21,14,11,
68,126,6,2,1,2,4,2,2,7,7,3,11,4,1,1,4,8,17,21,10,23,12,19,11,26,27,3,14,7,5,2,6,3,6,2,7,4,4,4,15,13,2,3,5,1,4,3,4,8,11,10,8,3,3,4,10,2,1,2,6,5,30,14,65,21,25,60,49,29,3,4,12,15,12,13,65,85,86,83,81,66,15,75,81,81,84,84,84,84,84,85,85,82,155,168,11,21,47,46,15,35,28,43,14,153,140,104,160,173,171,170,178,175,178,175,183,171,180,172,174,181,104,79,79,77,77,157,125,34,32,21,25,30,33,27,30,38,66,60,139,153,94,113,95,97,89,89,98,102,176,183,184,188,182,179,181,180,181,171,179,175,243,213,41,14,44,27,50,81,58,58,37,225,146,121,177,179,181,181,182,177,177,177,180,178,178,177,92,70,89,76,190,220,60,49,53,62,55,45,58,64,46,47,47,48,48,49,51,50,52,51,49,50,49,50,48,50,51,51,50,48,51,51,52,52,52,53,51,52,49,49,50,49,49,48,50,49,47,39,33,34,42,47,41,42,51,44,17,9,14,16,16,7,14,14,
120,108,5,9,2,3,2,3,4,3,9,6,3,5,5,4,4,6,31,93,10,33,38,19,15,19,34,22,12,6,10,3,5,5,10,7,4,4,7,4,11,6,3,2,7,3,3,2,6,2,8,9,1,8,2,3,1,0,1,3,2,2,9,15,16,15,21,13,15,10,14,6,10,8,8,4,11,83,85,83,80,68,16,76,82,84,84,87,85,85,84,86,85,84,146,160,19,29,46,50,15,57,31,51,16,127,157,94,112,159,160,151,176,177,178,181,179,177,179,173,177,178,103,83,78,75,98,72,77,39,32,20,25,28,29,25,33,36,60,56,92,87,191,145,107,109,108,112,101,183,180,184,182,183,185,180,180,179,182,177,178,178,247,216,38,14,35,30,53,67,54,50,24,223,121,113,180,178,182,183,182,174,178,180,180,179,180,179,88,71,90,77,181,230,67,80,15,14,41,83,54,52,64,61,47,43,44,41,46,47,49,46,49,48,45,44,45,44,46,45,46,46,47,46,48,49,53,50,51,49,49,45,47,49,51,48,48,50,49,47,46,41,37,30,32,42,45,42,47,52,46,51,51,54,52,54,
127,37,20,18,2,7,2,1,5,8,8,7,15,5,0,3,1,34,5,59,24,39,12,10,16,37,18,14,9,21,9,2,6,3,8,3,2,4,6,5,4,2,2,5,2,1,2,4,8,7,7,8,5,4,3,0,0,1,1,2,3,4,7,12,13,22,15,12,15,8,9,8,8,9,6,5,13,83,85,84,80,68,16,75,82,83,85,86,84,85,85,85,84,79,80,108,15,49,54,52,15,86,38,148,11,84,97,80,114,109,153,132,144,175,178,179,181,174,182,178,174,173,103,85,75,73,192,124,104,31,31,22,25,22,31,23,33,37,49,51,88,100,152,99,111,123,122,121,117,186,180,185,180,186,186,182,180,184,178,178,178,192,168,186,27,17,28,22,21,30,52,53,32,180,157,96,183,175,180,180,181,179,182,181,178,178,182,180,96,69,90,74,227,228,63,62,11,28,94,63,59,60,56,49,53,47,49,41,40,42,43,44,43,42,44,47,50,48,45,45,46,43,43,43,44,45,47,46,48,49,36,50,50,48,48,47,48,49,47,46,49,50,44,44,43,32,24,40,43,56,45,53,53,46,51,58,
126,64,9,27,2,2,3,2,3,4,7,9,8,4,2,2,1,5,7,30,48,38,32,44,15,10,24,15,10,18,6,4,7,22,3,5,9,3,5,6,12,5,3,3,5,6,1,4,6,4,4,9,5,5,3,0,3,1,3,5,6,10,21,9,22,15,13,9,15,7,8,9,6,7,4,9,27,88,85,89,83,70,16,73,81,82,85,84,82,85,83,85,83,80,81,109,6,13,13,14,14,28,43,31,10,86,82,75,81,139,129,137,119,154,178,181,180,180,181,174,172,174,112,75,64,60,153,173,88,24,26,20,24,23,26,23,32,35,50,43,91,95,179,144,103,106,109,107,76,182,183,183,176,182,184,182,184,182,180,179,180,187,181,161,53,46,59,80,41,125,59,67,33,167,183,95,184,177,177,185,183,180,181,178,176,178,182,182,88,72,91,71,213,227,11,18,8,34,43,40,45,23,51,48,39,49,58,47,47,42,43,38,40,40,41,42,42,43,44,44,40,38,41,40,40,41,39,38,40,42,44,46,47,44,45,45,36,50,48,47,48,48,48,49,47,45,42,38,27,26,39,40,38,46,51,50,
120,70,14,27,6,2,2,6,2,5,5,11,13,2,2,2,3,2,8,134,36,28,50,54,16,28,16,7,15,13,8,16,3,4,7,4,9,2,5,6,7,4,2,2,2,2,3,2,3,5,7,7,8,3,2,2,1,2,4,2,7,5,9,17,15,12,11,9,10,7,6,8,3,5,9,20,48,96,94,85,83,73,16,73,80,82,87,82,83,81,83,83,82,80,79,128,8,8,9,10,12,46,46,56,10,85,79,72,82,117,135,127,133,112,160,175,183,185,182,174,137,133,87,68,46,38,73,82,67,27,24,23,18,26,27,25,28,31,34,48,154,162,106,102,100,91,91,101,108,138,186,181,176,183,184,184,179,178,181,177,172,192,163,179,22,25,24,29,24,26,25,27,31,178,106,96,180,179,178,182,180,179,180,177,178,182,182,180,84,74,91,75,227,60,8,16,15,29,34,47,23,23,14,46,50,43,38,50,58,51,50,40,39,38,40,43,42,41,45,44,45,47,45,46,45,45,45,42,43,42,42,43,46,45,46,45,47,45,75,46,45,46,48,47,51,49,49,47,45,43,39,23,23,37,42,38,
120,103,33,21,3,1,2,6,1,7,5,7,2,2,2,2,1,2,5,34,34,37,52,41,36,34,24,12,10,7,7,11,7,8,5,5,2,6,2,4,2,2,2,2,2,2,3,1,2,2,5,7,2,4,7,0,1,3,4,4,3,10,15,12,13,10,16,11,7,11,8,4,5,6,14,15,45,115,116,104,91,73,23,73,79,82,82,82,81,81,82,81,78,84,118,111,85,90,95,112,119,129,126,85,82,111,120,84,84,89,111,116,124,122,106,153,178,183,182,178,21,20,17,17,15,17,17,16,14,18,30,23,26,20,21,23,24,24,51,50,149,154,100,108,112,111,111,111,112,103,185,179,181,186,185,182,177,181,185,182,174,206,185,196,58,74,88,96,111,113,114,117,112,192,166,100,181,180,182,181,179,180,180,181,178,180,177,178,83,77,95,77,197,222,11,6,9,14,10,14,11,8,15,43,33,41,49,41,40,50,53,41,46,36,37,37,37,38,41,42,45,42,44,47,43,42,43,42,45,43,40,40,42,44,44,46,47,51,28,42,43,45,46,46,47,48,49,48,50,50,46,44,40,34,25,37,
97,94,54,49,6,3,2,3,3,6,3,8,3,4,2,3,3,3,14,23,19,31,35,21,26,17,19,9,9,9,11,7,6,8,2,4,3,6,2,3,5,1,2,0,3,2,2,3,2,3,8,5,7,4,6,6,3,1,7,6,5,5,12,9,17,10,4,8,15,6,4,3,5,17,19,20,48,102,122,124,96,91,20,72,78,81,81,75,81,80,80,80,75,144,144,145,142,139,144,139,141,142,138,144,139,145,148,137,78,84,89,102,106,112,113,101,140,167,187,176,13,19,19,18,17,17,16,18,15,18,29,25,36,24,35,29,32,36,54,47,148,153,100,182,105,106,105,100,98,170,183,178,182,188,182,182,177,183,181,183,183,226,229,226,227,223,216,225,218,222,214,225,223,223,222,220,171,181,179,180,181,181,180,180,180,178,174,178,87,79,94,77,200,219,26,9,4,13,10,9,6,8,17,33,19,13,38,49,49,39,37,48,55,44,46,34,36,37,37,40,38,41,44,44,41,43,42,44,44,45,41,41,40,40,40,41,51,195,129,56,46,47,48,49,49,48,49,51,50,50,50,50,49,47,47,46,
141,67,59,59,13,1,1,2,1,5,6,6,3,5,5,4,1,4,6,8,16,17,21,16,14,18,9,7,7,5,10,6,4,5,5,5,3,6,5,2,2,1,1,1,0,2,3,2,2,5,16,4,1,9,7,6,2,6,5,3,9,8,8,11,12,11,8,12,9,4,2,11,18,17,19,19,83,89,110,143,116,85,17,71,78,79,79,76,79,79,79,79,78,107,108,104,100,95,96,102,92,97,91,103,104,107,118,105,78,80,86,86,95,97,98,120,113,139,157,174,16,26,12,21,18,22,18,19,19,22,31,25,30,50,28,31,33,37,54,49,150,155,102,181,120,113,107,122,117,175,184,181,183,182,181,185,185,182,179,183,182,229,224,220,222,224,225,221,220,220,223,230,222,220,227,216,102,146,178,184,183,182,179,179,181,181,175,177,76,77,93,76,229,204,61,8,7,3,10,8,9,11,14,12,24,14,31,38,39,50,51,38,39,53,51,44,52,36,38,34,35,45,72,41,40,40,42,42,42,42,43,45,46,42,43,41,149,165,109,85,133,168,201,200,197,199,206,205,206,209,216,219,216,217,218,217,
142,92,75,69,10,3,2,2,1,2,3,2,1,0,0,0,0,0,0,1,2,6,4,11,17,8,7,7,0,4,7,6,9,4,2,2,3,2,2,2,2,1,1,3,1,1,6,2,1,5,6,7,3,7,8,3,4,7,13,9,15,11,11,8,8,16,6,11,3,7,13,18,23,23,22,22,52,137,114,108,147,103,18,70,76,77,80,77,77,76,77,76,77,76,76,75,74,75,77,75,78,85,84,78,75,75,76,77,81,80,82,86,82,88,95,99,117,138,128,135,156,163,107,63,63,55,56,95,112,29,29,22,30,24,27,26,29,36,45,48,148,159,104,169,104,103,118,114,92,183,182,182,178,177,183,185,185,178,181,183,182,177,105,108,105,101,104,103,101,102,105,104,104,106,104,101,102,105,183,179,182,182,177,180,181,184,175,177,78,75,92,77,49,229,73,7,6,2,5,3,6,8,10,9,17,6,19,49,42,39,40,49,48,37,38,53,52,48,50,33,38,35,99,41,37,42,41,42,45,42,43,43,42,46,43,46,110,127,114,113,81,91,97,110,117,126,131,143,153,161,172,183,186,194,202,210,
139,122,77,60,26,5,3,3,2,2,3,0,0,5,4,3,2,7,15,8,2,1,0,1,4,5,6,4,9,8,8,6,8,1,1,2,3,8,3,4,2,1,2,0,3,3,1,1,2,6,6,3,2,8,4,6,6,11,10,12,16,12,8,21,8,13,11,8,5,13,29,30,26,26,24,25,49,101,134,134,89,122,20,68,74,75,139,89,77,76,75,76,76,76,76,76,76,76,78,77,77,84,84,76,77,76,78,77,78,78,83,81,88,80,86,102,96,102,109,98,112,134,98,72,71,65,60,106,125,28,20,21,29,22,22,25,26,31,35,45,150,158,98,109,84,76,76,101,111,136,177,182,181,183,185,186,182,180,180,183,179,175,180,118,111,109,106,106,106,105,106,106,109,107,107,107,103,104,184,180,177,181,178,179,180,182,176,177,82,75,95,81,223,160,41,11,6,8,5,1,2,9,6,12,17,11,6,38,42,50,43,39,49,44,43,36,43,53,47,40,37,34,139,34,32,39,42,47,44,42,43,43,41,40,43,39,132,124,107,107,42,46,46,46,48,50,49,45,42,42,45,43,42,43,44,42,
139,116,72,54,41,4,1,1,1,2,2,1,4,7,2,5,3,2,6,19,15,7,7,8,2,1,2,0,2,8,7,8,8,4,4,4,5,4,2,2,1,1,4,5,4,1,2,3,5,1,2,2,3,6,5,3,9,9,8,14,17,13,10,6,14,8,10,9,13,28,27,25,22,22,24,23,52,86,100,122,132,95,17,66,73,73,77,109,94,75,75,74,75,76,75,76,75,75,75,76,77,80,81,76,77,76,78,77,77,77,82,79,79,87,81,87,101,94,87,90,79,89,61,74,73,67,63,109,124,29,27,18,25,25,29,25,27,33,48,45,151,160,98,112,115,106,110,118,108,102,184,182,183,178,183,186,183,180,184,180,181,182,180,183,181,185,182,181,182,183,180,182,185,185,185,186,181,181,180,182,179,184,178,180,183,177,180,180,91,74,96,81,201,220,28,23,18,13,8,3,1,3,6,5,16,14,12,21,24,41,46,45,37,35,48,46,39,37,50,49,46,42,107,31,33,34,34,36,39,41,39,42,41,42,42,42,111,118,107,106,43,39,42,42,44,45,45,46,47,42,42,43,42,42,43,44,
119,111,75,9,3,5,2,1,1,2,4,3,3,4,4,3,5,0,6,12,14,4,5,9,8,5,3,0,2,2,8,1,0,2,4,3,4,3,1,4,2,4,4,3,3,5,2,1,2,1,4,6,5,4,4,9,6,15,13,14,9,10,9,11,11,4,5,13,29,33,29,27,24,23,21,25,51,80,86,109,129,103,18,65,71,72,80,78,130,86,73,73,74,73,73,77,74,74,75,74,74,77,77,74,75,75,76,77,76,78,76,80,79,79,82,82,88,93,85,75,79,72,46,82,70,69,61,108,122,32,28,20,24,22,29,21,27,27,48,43,153,161,101,157,113,115,115,116,102,166,186,184,182,179,181,184,183,182,182,183,179,178,181,181,183,182,177,181,182,182,183,183,183,184,183,184,180,179,177,183,180,183,180,181,179,178,177,181,100,75,96,82,217,215,32,28,22,21,15,8,7,5,11,4,30,16,12,8,11,16,23,48,44,43,35,40,48,49,39,37,43,48,123,40,33,26,32,35,31,36,38,41,43,43,43,41,124,116,131,109,42,42,42,43,44,44,43,44,43,44,44,42,42,43,41,40,
41,2,3,10,53,20,2,1,2,1,3,7,4,4,4,4,4,1,3,4,8,5,6,6,7,5,8,3,1,4,4,8,5,4,2,4,3,2,0,2,4,3,3,7,3,4,2,4,2,2,2,3,4,3,6,9,13,14,22,10,10,9,9,10,13,15,14,28,35,34,34,25,26,27,25,22,56,80,78,80,97,132,20,63,70,70,87,86,80,120,90,71,72,75,73,72,76,74,73,72,77,72,73,72,73,73,74,73,75,75,75,75,81,80,80,83,84,88,83,70,62,67,33,67,64,59,152,145,114,36,24,17,22,21,28,20,24,22,40,41,154,159,103,173,169,104,103,107,107,181,186,183,183,181,183,183,183,183,183,186,182,181,182,180,181,178,181,181,183,183,182,185,186,184,184,187,183,181,181,183,183,182,179,182,181,174,182,184,111,74,96,79,221,227,27,31,33,32,30,21,15,4,11,10,11,19,20,7,17,9,17,35,33,37,37,39,35,42,49,48,38,41,142,47,41,39,33,31,34,36,35,36,39,43,40,41,108,117,108,105,38,39,40,40,40,44,41,40,41,42,45,41,44,42,43,43,
40,58,66,63,28,11,8,0,1,2,3,4,6,6,6,6,4,8,5,9,6,7,5,4,3,6,2,7,0,2,5,4,6,7,6,7,2,1,3,1,2,3,5,1,2,4,3,2,3,2,2,2,2,1,4,6,12,14,21,9,11,10,10,6,6,28,40,35,44,37,21,26,27,26,26,22,57,77,77,75,75,70,22,62,67,69,92,80,95,85,83,93,75,70,74,70,68,71,70,69,65,70,68,70,70,70,71,70,72,72,72,72,72,80,79,80,87,84,87,74,60,43,25,41,38,41,82,92,81,34,24,16,22,23,27,20,25,19,40,41,151,159,101,173,182,179,181,178,183,177,180,185,186,175,181,186,185,180,181,184,182,182,183,181,181,175,177,181,177,179,181,184,182,187,185,184,185,181,178,184,183,180,185,184,184,180,184,184,124,72,95,81,223,180,25,23,25,26,30,30,23,23,11,14,20,5,22,12,10,11,27,29,42,39,34,53,51,52,49,54,48,46,149,44,50,50,53,40,33,33,38,40,37,37,39,39,121,120,106,105,44,41,44,40,39,43,46,48,47,47,56,66,69,73,61,63,
105,59,60,38,26,27,8,2,4,2,2,5,8,10,6,4,5,14,2,6,6,7,6,5,4,1,1,2,1,2,4,2,2,5,8,4,3,3,3,2,0,2,0,2,3,3,6,4,3,5,3,1,1,0,2,9,7,16,13,5,10,10,4,9,29,38,34,24,32,33,30,24,23,26,19,23,94,89,76,75,73,65,14,60,65,66,84,93,106,94,82,72,81,78,68,76,71,67,68,70,63,64,67,68,69,68,69,67,69,70,71,71,72,72,78,78,80,87,76,72,66,58,38,58,59,50,53,107,101,29,22,17,24,26,27,22,27,28,36,40,154,158,106,160,182,180,177,181,185,181,179,185,194,172,180,183,178,176,181,186,182,183,186,181,177,177,180,177,174,178,179,178,184,187,186,188,186,178,176,179,183,183,184,187,179,179,180,178,143,54,95,84,206,227,28,27,33,32,30,28,31,29,27,14,10,8,17,7,8,11,17,20,33,113,121,42,42,37,41,45,52,49,159,44,40,42,48,48,42,51,29,32,35,39,38,37,113,121,109,103,42,41,43,44,43,43,43,45,47,43,43,45,45,45,45,48,
119,67,59,31,40,27,2,3,3,9,6,4,13,17,8,6,5,6,3,7,14,5,4,13,0,3,8,2,1,3,5,4,5,2,2,2,2,2,2,2,3,5,1,2,3,7,6,1,3,5,1,3,1,1,1,8,10,17,16,12,8,7,8,27,34,30,28,31,33,26,23,22,25,25,25,30,62,128,104,70,68,61,11,56,58,63,76,93,97,112,74,84,71,73,82,67,75,69,64,67,68,63,63,66,66,66,67,67,67,67,68,69,72,72,70,72,72,76,76,71,68,65,46,61,58,51,45,86,103,33,23,17,25,26,26,21,26,33,35,44,158,163,106,139,184,182,185,183,183,184,184,181,184,180,187,186,183,182,186,186,187,187,186,184,177,167,174,175,165,177,176,175,186,190,186,184,183,181,178,186,191,184,188,182,182,182,181,183,151,66,97,83,190,223,31,26,32,31,31,31,30,31,30,27,24,23,10,9,14,19,18,12,40,88,65,49,43,44,50,51,47,46,162,51,55,45,44,49,53,49,49,48,34,33,36,37,113,121,110,109,44,44,44,45,43,46,44,46,43,44,44,42,43,45,44,45,
83,68,71,51,38,13,0,0,3,3,10,11,14,12,10,6,6,12,21,12,8,9,12,21,3,3,4,4,3,2,4,2,0,1,1,1,2,2,5,2,6,6,1,1,4,6,3,4,2,1,2,1,0,4,3,8,28,40,19,28,4,7,21,34,35,36,34,29,32,34,30,29,24,22,34,33,70,74,141,116,63,51,11,47,56,56,95,80,97,107,111,74,81,66,70,88,65,70,64,61,61,64,61,62,62,61,62,65,64,65,64,66,68,72,67,66,68,68,76,70,70,61,39,63,55,53,49,92,94,29,21,15,24,24,26,20,26,32,30,46,158,164,104,162,186,188,195,187,187,191,187,191,189,190,194,191,192,201,189,191,194,196,198,197,180,137,160,173,171,175,179,149,189,203,188,188,173,189,184,190,181,204,195,191,191,193,183,182,155,64,93,81,226,232,29,33,30,30,33,34,34,40,38,32,24,22,15,10,10,9,53,73,148,188,80,85,107,95,113,138,157,180,165,200,202,197,195,200,201,201,199,210,206,127,48,32,120,118,110,110,46,47,47,46,45,45,43,45,45,43,45,44,43,46,45,46,
92,81,55,53,66,1,1,3,7,9,8,7,5,5,7,11,6,25,24,5,12,30,14,12,10,9,5,3,5,6,2,2,2,1,1,1,1,2,2,2,4,3,8,6,3,2,2,2,0,1,0,1,1,3,4,31,36,33,51,8,11,39,43,42,35,33,30,35,31,27,33,37,24,23,25,28,134,107,85,51,97,61,10,49,53,52,100,93,71,83,88,76,62,60,62,56,81,64,81,61,63,64,72,74,64,57,57,57,58,59,61,60,62,62,67,64,54,56,58,81,68,62,33,49,47,50,57,62,70,21,17,14,21,18,20,19,23,29,39,52,130,122,113,208,212,214,222,202,200,204,172,215,186,207,199,200,207,183,214,206,203,197,244,229,225,174,187,188,180,177,174,182,184,231,229,159,220,221,184,200,159,208,166,205,203,196,193,190,163,55,57,70,123,224,25,35,32,33,28,33,33,38,34,37,29,29,24,23,6,23,49,123,74,53,134,176,130,111,199,204,211,222,179,127,158,181,197,201,197,203,209,206,208,203,215,90,116,120,108,110,66,86,86,101,90,53,77,89,86,62,63,101,109,135,189,191,
1,3,29,65,52,1,0,2,15,10,16,28,10,9,17,14,11,6,2,14,24,39,20,13,3,9,6,2,3,3,2,1,1,0,1,1,2,2,1,2,2,3,4,4,4,2,2,1,1,1,2,7,5,3,10,46,68,40,67,13,33,42,45,37,32,35,36,37,31,30,44,45,47,48,37,31,86,69,59,52,66,102,10,47,47,45,67,64,70,55,46,51,72,61,58,65,54,54,53,48,42,43,48,48,59,60,54,46,45,51,50,50,50,60,55,52,53,53,52,46,58,47,29,44,46,121,44,82,40,19,13,13,18,15,16,19,19,26,33,50,83,88,141,210,197,139,202,168,161,115,154,159,139,161,188,196,182,188,217,169,187,166,250,147,107,110,111,106,111,112,114,107,103,104,102,95,91,158,188,143,212,176,176,155,192,199,186,146,209,48,91,136,113,123,21,39,41,42,41,43,46,40,41,38,37,37,39,35,26,57,151,111,156,157,226,210,205,202,202,202,204,208,212,209,206,202,202,199,196,198,204,107,207,216,222,219,126,118,106,111,187,189,197,198,199,196,198,180,144,131,140,159,168,175,178,184,
3,0,0,1,1,1,0,10,15,9,10,24,24,10,9,7,3,7,8,11,7,18,8,16,17,9,6,3,2,4,2,2,0,1,1,1,2,2,1,3,6,5,3,4,5,1,1,2,1,3,1,3,7,15,6,19,16,19,14,40,50,50,38,38,39,46,44,43,46,68,107,102,144,131,136,172,83,58,69,56,81,44,8,41,39,37,46,37,41,43,42,44,49,55,47,64,82,59,55,37,47,51,49,49,42,53,44,48,45,32,37,43,43,49,45,40,55,43,52,50,33,30,23,40,42,62,60,75,38,24,21,24,22,19,12,17,19,27,41,65,77,86,156,174,98,172,133,132,113,127,188,117,194,156,171,173,133,200,213,171,178,198,242,237,126,103,107,107,105,106,101,98,99,92,109,77,55,65,192,159,196,205,128,175,186,157,181,93,172,63,84,76,60,115,23,40,47,45,47,52,51,49,54,50,51,52,54,54,46,117,159,214,111,111,224,205,206,200,209,204,203,199,202,204,192,186,181,174,162,153,141,44,142,154,168,168,175,144,121,131,157,97,79,76,98,116,137,146,150,155,158,171,188,187,186,186,
78,72,8,0,0,1,0,5,14,10,11,20,41,8,8,15,32,41,25,39,42,22,0,10,7,5,4,2,1,4,2,2,0,1,0,1,4,0,3,1,4,5,6,0,2,0,3,1,0,2,1,2,6,26,10,10,14,16,47,122,178,164,188,195,190,188,190,188,171,163,183,182,195,192,179,189,61,74,52,33,53,52,8,37,40,35,48,60,42,34,55,47,49,47,60,46,61,66,64,51,87,61,50,48,42,40,47,42,53,47,36,39,45,42,43,46,56,56,53,63,33,46,35,39,33,53,44,96,37,8,32,30,34,47,53,59,63,68,80,70,89,102,179,143,224,211,220,227,93,104,80,98,157,111,144,148,137,173,146,147,181,189,227,241,159,186,160,185,174,178,178,178,112,191,165,104,61,61,75,193,218,216,221,213,191,199,215,159,166,54,48,50,122,206,183,218,216,210,211,221,219,39,210,218,223,220,218,218,213,218,199,201,128,205,126,168,135,48,38,55,118,78,49,44,46,102,64,152,180,206,200,57,202,203,206,198,191,191,165,174,164,191,190,194,198,199,199,198,194,194,193,192,189,188,186,187,
100,18,5,1,1,1,3,16,13,3,18,6,2,8,17,35,36,20,51,47,34,41,40,44,12,3,2,0,5,2,2,1,2,0,3,1,2,6,2,0,4,4,3,1,2,6,6,1,1,2,1,54,13,15,56,171,158,183,185,185,200,198,193,203,196,181,164,190,180,197,200,205,150,151,135,108,38,40,47,71,40,60,7,38,32,28,33,47,51,46,38,37,39,35,39,29,65,89,105,43,97,112,78,47,31,27,49,65,37,56,48,40,40,40,32,33,34,44,48,80,75,50,28,28,42,47,41,81,47,50,75,64,57,108,165,184,152,142,137,148,207,215,213,108,174,125,144,102,169,192,170,186,194,203,211,226,215,221,227,224,219,229,243,228,133,168,143,152,156,157,171,163,142,155,141,126,60,66,72,82,237,211,231,239,237,233,237,235,227,230,228,177,221,212,221,208,209,215,226,222,201,42,220,202,224,221,216,216,215,223,224,207,202,155,43,42,40,180,42,43,49,52,182,50,47,46,47,125,99,180,199,96,207,192,200,200,192,196,192,206,170,176,182,175,187,193,195,198,197,201,196,187,166,152,174,193,
77,2,15,0,2,1,4,59,39,5,10,25,78,78,135,179,91,90,199,174,175,189,171,159,168,145,22,9,9,6,3,1,1,1,0,5,4,1,1,2,7,1,3,8,3,2,0,1,0,1,5,2,2,56,108,131,166,168,172,164,168,180,175,171,172,184,194,190,202,202,201,209,173,212,190,208,148,92,101,94,84,52,68,22,58,52,54,51,52,56,52,46,52,50,66,68,53,54,49,58,57,53,58,61,61,50,52,55,66,90,81,65,92,122,111,70,86,118,186,168,129,71,77,49,123,114,85,82,93,102,125,164,147,149,149,167,190,195,214,218,216,222,227,94,221,224,234,220,224,226,232,216,229,231,229,215,227,228,222,217,229,214,228,181,193,197,211,218,213,230,224,228,228,232,235,215,226,195,212,225,233,226,226,233,228,226,228,236,233,235,227,170,207,218,217,218,217,215,208,217,225,38,222,227,229,217,213,210,205,216,211,173,83,190,145,91,89,153,45,174,190,199,200,196,191,203,199,208,208,207,205,49,200,203,200,201,177,190,192,63,167,184,189,195,184,189,195,194,190,191,191,189,189,189,182,164,
14,66,3,1,1,3,1,6,4,115,146,109,54,30,113,65,89,144,155,193,195,177,180,193,197,196,106,11,24,7,4,1,5,2,3,3,5,4,6,2,2,6,2,6,3,3,0,1,1,0,2,12,7,62,38,115,157,163,164,169,150,152,167,166,175,174,196,190,192,196,198,203,195,195,163,122,89,113,107,178,175,127,113,23,123,122,88,64,41,45,70,90,88,120,104,57,67,61,68,67,65,70,85,78,82,73,79,58,60,82,114,119,125,143,152,156,164,175,171,115,84,95,117,49,159,167,187,205,194,212,211,213,217,212,213,210,207,206,215,216,216,209,219,133,220,229,218,225,226,228,227,220,218,214,229,229,229,226,231,221,221,211,225,220,222,222,226,227,225,187,209,220,225,226,224,225,203,220,225,227,228,229,203,230,219,215,218,221,225,233,228,36,40,222,218,218,218,220,222,214,216,113,194,179,173,125,81,125,183,188,182,185,185,194,194,191,200,195,103,191,190,198,198,199,197,195,191,211,211,213,212,62,211,204,198,200,200,197,194,104,33,166,178,142,184,188,191,169,195,192,189,188,187,188,185,183,
7,21,2,1,1,4,2,7,88,146,181,160,128,25,32,94,90,182,178,158,186,191,200,192,187,157,108,14,22,6,4,1,3,1,2,7,2,5,6,4,7,11,2,5,3,0,1,1,1,1,0,1,7,68,49,88,169,165,162,160,169,171,172,174,179,173,174,170,150,169,164,157,142,135,104,129,99,114,126,137,144,120,113,25,107,88,51,62,109,166,201,206,200,174,130,89,58,56,57,78,64,62,75,96,93,79,72,88,59,69,108,103,117,153,207,215,207,211,210,210,210,207,206,102,214,211,217,214,212,213,206,208,212,204,215,207,201,207,210,212,208,213,219,164,217,221,221,226,217,219,220,220,222,220,223,230,233,229,232,232,220,203,224,212,224,226,220,217,220,227,222,186,218,219,206,216,218,218,225,224,225,229,207,228,228,226,217,201,213,179,174,83,79,94,130,186,204,203,133,157,192,46,188,186,186,188,188,196,195,199,196,193,193,196,196,195,194,199,98,200,194,194,202,194,193,196,194,194,195,184,168,62,182,173,195,201,196,190,186,60,29,35,181,189,196,187,180,186,179,193,188,185,185,187,185,184,
11,5,4,2,4,2,14,7,78,166,187,195,203,90,115,155,178,179,205,204,209,189,190,187,169,162,199,10,28,5,6,5,5,8,5,5,3,4,8,7,10,13,8,3,5,4,1,1,3,1,3,6,11,37,36,78,68,83,57,75,102,138,159,146,159,188,171,185,188,187,180,185,185,198,216,210,201,212,219,222,215,193,186,68,216,210,191,190,171,194,192,199,169,99,108,125,128,119,142,151,142,149,181,57,61,53,65,62,93,167,201,214,207,209,215,209,211,208,210,208,212,203,206,85,212,213,208,195,208,208,205,198,172,169,147,130,123,128,147,177,197,200,140,109,203,203,205,201,202,203,205,205,208,204,205,207,206,203,203,202,201,195,209,207,216,219,212,212,209,205,205,200,202,209,205,207,205,204,204,196,197,198,201,199,196,199,196,194,201,201,199,199,196,180,171,196,193,196,191,195,132,46,196,193,194,193,201,202,203,196,190,194,192,191,192,191,193,190,74,197,199,192,190,191,192,190,196,193,191,189,186,92,193,191,191,177,190,186,180,54,37,33,186,187,186,188,186,186,186,190,190,189,187,186,185,187,
3,2,0,1,7,14,9,53,140,167,176,175,180,158,189,181,132,174,176,175,177,174,169,174,158,148,116,5,8,9,5,3,6,7,9,27,6,5,12,10,7,6,6,20,7,5,1,2,5,13,15,9,9,98,66,107,180,178,184,184,181,186,192,190,185,191,187,188,186,189,190,190,195,194,195,192,191,187,187,186,191,187,187,23,182,190,189,190,192,192,196,192,196,192,190,197,194,193,192,194,200,192,187,187,183,152,189,191,193,177,191,189,188,190,190,194,195,187,141,97,92,86,66,42,117,161,170,176,193,199,200,204,202,196,198,199,199,197,203,120,205,204,204,84,205,207,122,204,204,207,204,208,205,206,209,202,206,209,207,206,207,193,209,209,205,204,205,202,205,203,204,203,205,206,204,202,202,198,199,201,202,199,199,203,201,199,203,204,204,204,204,201,194,191,131,201,192,192,189,194,193,30,203,198,193,191,190,193,189,190,192,192,193,188,190,188,192,190,68,186,189,188,189,188,190,189,188,191,189,189,192,125,194,192,193,214,192,193,49,43,20,70,186,189,191,180,178,170,181,185,187,191,193,193,198,184,
2,0,2,1,10,196,202,82,198,179,202,202,101,159,172,207,203,206,202,197,198,204,200,189,159,79,32,13,12,7,5,61,6,6,14,5,10,10,28,17,12,14,36,14,10,3,3,49,8,55,84,111,11,113,47,189,198,201,202,200,202,200,204,203,205,201,206,203,203,206,202,198,202,206,207,207,203,182,205,205,203,206,205,20,172,204,205,208,210,211,129,194,210,210,210,206,212,205,206,217,216,211,210,178,155,83,66,59,58,65,96,149,187,192,197,199,201,202,195,192,194,191,194,71,193,196,196,195,198,195,191,190,194,194,196,194,177,177,200,103,194,195,195,84,194,196,112,197,201,201,194,197,197,199,199,199,194,199,197,199,199,176,202,200,200,198,200,200,198,200,198,197,197,197,198,198,200,199,198,200,198,202,186,194,196,197,196,195,193,195,196,194,195,193,192,129,192,192,193,190,193,36,116,194,190,191,188,188,195,184,183,190,191,186,183,190,189,193,71,188,188,191,188,194,190,187,189,188,185,183,182,70,193,194,154,195,192,190,41,34,36,176,182,187,188,186,176,168,180,183,179,180,181,177,181,182,
1,1,1,2,29,101,169,62,158,173,162,164,121,139,176,176,178,176,179,180,153,179,176,165,137,128,19,8,8,6,5,1,2,10,29,124,179,75,35,13,6,9,4,1,4,71,21,9,16,45,167,172,35,81,125,180,186,189,189,189,191,193,189,191,195,195,197,196,196,199,196,197,195,201,198,201,197,201,201,202,192,199,201,21,195,193,194,197,197,199,109,206,204,205,201,202,206,206,204,211,205,207,211,214,210,44,210,202,201,200,205,208,201,205,199,201,203,202,202,203,198,199,201,38,203,201,201,200,203,201,196,202,197,196,199,201,199,197,202,103,195,199,201,151,201,204,136,161,203,202,202,200,202,190,202,200,202,200,200,198,194,135,200,197,197,195,198,198,198,198,200,199,198,194,197,193,197,199,197,202,204,208,122,202,201,198,202,199,195,195,195,193,196,198,196,197,136,188,188,190,187,59,189,120,197,189,190,192,195,186,190,191,191,190,187,192,186,190,179,190,191,196,199,195,188,193,193,190,192,186,185,68,186,97,196,185,198,84,76,49,172,181,184,192,193,188,195,185,187,182,191,176,139,153,149,194,
0,1,1,44,125,97,154,93,175,197,196,182,156,192,183,182,189,155,78,21,6,7,7,7,8,8,4,0,4,4,4,60,46,81,107,170,176,120,41,45,136,42,37,81,36,11,8,26,108,162,157,155,37,197,190,173,192,191,201,195,192,194,192,190,201,197,200,199,199,198,199,201,199,200,194,196,192,193,196,195,197,196,112,45,190,196,198,199,197,119,155,193,199,198,198,192,188,189,190,185,196,196,195,193,195,67,193,192,191,196,195,194,197,197,195,199,199,201,194,191,190,191,187,55,190,191,191,188,191,189,181,194,194,195,196,194,193,198,197,169,122,200,193,65,196,200,201,110,199,202,200,197,198,197,198,201,200,199,197,200,199,155,199,199,201,199,197,198,198,195,196,197,195,197,196,197,198,199,196,198,200,194,193,200,200,195,196,197,197,195,196,198,198,197,193,192,189,136,194,192,189,35,195,189,123,190,188,189,187,183,186,189,192,192,188,187,189,186,83,193,191,194,193,201,202,196,194,193,187,195,192,80,196,196,194,182,71,152,166,201,180,113,192,189,190,187,187,183,169,172,176,111,158,180,171,139,
0,0,3,2,2,20,103,95,140,180,181,176,143,137,94,23,9,10,8,10,10,144,163,172,108,161,175,6,8,10,8,46,68,155,179,185,195,206,148,86,104,55,42,59,125,163,188,115,145,130,167,178,35,173,183,183,185,181,186,185,179,190,191,193,189,193,185,196,194,195,194,199,189,187,192,190,192,196,194,197,198,200,95,36,195,195,195,196,204,111,200,196,198,199,198,201,195,196,196,196,197,198,191,195,194,125,194,195,181,199,199,198,200,197,198,198,197,197,195,194,197,197,195,67,193,195,197,197,196,195,196,197,197,192,195,197,195,198,197,191,104,203,200,76,196,200,199,104,200,202,201,199,202,197,197,201,204,204,202,203,196,125,201,199,201,202,201,205,204,202,202,202,201,199,200,199,196,201,200,203,199,198,173,198,198,199,199,199,200,207,207,206,206,204,206,203,201,199,121,189,188,41,187,183,187,109,198,192,194,193,191,189,191,189,189,190,188,183,94,183,191,191,191,193,199,195,196,195,188,163,198,151,100,188,86,35,97,122,174,175,132,94,159,183,195,164,167,142,173,145,160,154,184,140,135,154,
0,1,6,7,3,2,6,12,63,70,128,113,80,27,5,10,114,112,96,64,38,186,134,99,147,190,166,44,36,25,7,37,16,121,166,161,192,184,191,102,117,38,91,70,90,179,149,192,189,191,191,188,33,191,185,188,185,190,190,191,191,192,184,194,194,193,192,191,193,193,195,192,194,195,197,200,198,197,196,194,193,99,198,37,198,197,197,197,145,146,192,195,192,198,200,202,198,197,202,200,197,199,198,199,198,103,191,190,192,193,191,187,191,191,191,192,191,194,202,202,200,200,199,59,201,204,204,204,202,203,199,201,203,200,203,201,203,199,202,202,126,204,202,83,197,202,205,130,169,203,203,201,200,202,201,202,203,201,205,205,204,76,204,200,204,203,204,205,207,204,204,203,205,206,208,206,206,206,205,204,204,187,72,204,204,203,205,206,206,204,204,207,203,200,177,175,199,201,200,147,193,52,195,194,190,187,130,190,187,197,196,194,194,191,190,195,194,194,133,191,192,190,192,193,181,187,188,187,187,184,188,135,61,106,138,166,151,88,151,151,195,193,195,128,192,193,189,197,198,197,197,197,184,173,166,150,
1,3,37,88,103,5,5,5,3,8,4,5,6,2,16,120,75,91,84,97,63,92,76,112,199,162,139,26,32,31,60,22,43,91,138,165,179,198,202,206,66,192,108,129,74,97,207,194,207,193,197,185,27,193,196,193,195,194,186,194,176,195,196,199,189,200,198,202,200,204,199,198,194,197,198,199,198,203,202,204,188,95,193,40,199,202,204,199,107,207,207,209,207,206,205,199,208,207,209,210,208,207,203,208,208,32,204,205,206,205,206,207,211,208,203,199,187,156,113,160,205,208,205,26,203,206,206,201,206,203,186,145,104,136,175,175,179,203,203,203,117,213,209,62,205,205,202,185,82,113,103,114,162,163,166,192,207,208,204,206,169,34,161,140,111,104,122,158,167,175,189,199,200,206,199,200,198,199,203,205,204,147,107,86,137,156,159,169,189,192,195,195,198,193,193,194,200,192,198,202,156,94,89,111,113,100,99,88,136,145,175,160,150,154,116,132,205,194,112,112,151,113,93,104,152,159,146,93,42,41,36,32,123,133,129,148,159,200,187,189,179,196,166,173,181,196,195,194,197,191,186,190,193,189,175,155,
3,18,11,15,111,36,147,5,78,136,156,32,66,56,66,60,88,107,106,114,75,45,94,170,197,177,82,15,63,4,82,33,45,65,78,194,185,111,99,126,177,49,82,157,151,207,207,193,207,206,206,207,15,208,186,207,204,206,192,153,116,102,93,123,177,189,192,205,209,210,208,209,209,205,212,210,205,206,204,193,127,172,182,50,154,162,165,118,53,115,166,180,187,193,196,189,195,191,195,195,195,197,191,191,157,57,130,176,181,187,191,193,197,163,203,197,197,195,198,194,191,191,179,89,152,197,198,192,192,191,197,198,197,197,197,196,193,193,195,196,193,198,194,187,193,200,197,198,198,195,196,172,195,196,194,192,184,189,181,182,193,187,89,182,182,178,177,179,177,184,182,188,180,149,184,176,181,173,147,179,176,182,181,177,169,170,174,169,168,161,161,165,174,165,170,167,163,162,161,157,141,164,166,168,172,168,211,188,185,193,190,193,190,192,190,193,189,174,156,152,148,131,135,85,57,51,44,37,52,70,129,140,153,192,193,195,198,192,196,173,195,185,186,174,199,187,174,174,190,191,189,191,190,183,176,185,
38,34,0,5,30,8,178,65,60,134,163,99,10,96,41,43,73,42,29,105,84,3,30,114,65,69,49,26,25,16,6,15,9,79,68,159,185,93,161,188,139,59,94,144,181,176,143,183,181,181,181,149,78,169,180,177,174,178,176,183,183,183,184,184,165,193,191,188,186,195,201,192,199,198,200,190,190,195,191,183,179,195,193,189,190,186,199,199,210,197,182,145,176,161,154,155,156,174,172,181,176,181,129,174,173,167,167,164,169,163,162,154,155,111,147,145,128,126,108,109,93,107,107,91,112,112,114,96,95,79,85,84,77,84,76,66,97,92,82,87,99,104,109,105,101,91,108,93,93,101,97,100,99,109,98,105,101,102,100,98,101,106,65,100,104,99,95,97,92,100,95,101,103,71,92,92,96,95,96,100,99,95,96,97,90,89,90,85,93,92,94,93,95,86,89,89,92,91,100,92,94,91,90,89,86,87,174,75,74,80,80,68,50,50,45,40,33,42,44,43,140,43,40,134,142,162,180,184,127,201,190,194,193,191,195,194,194,195,196,197,196,209,198,184,189,195,191,194,196,197,191,191,189,189,193,193,
35,43,1,5,13,15,129,137,19,110,157,108,12,20,20,28,8,14,33,82,107,49,2,38,50,31,142,60,49,58,8,18,9,7,77,92,25,83,26,50,11,77,114,90,117,94,117,97,103,113,116,113,96,112,126,134,126,128,68,97,107,104,99,88,102,108,115,112,118,103,102,116,122,114,121,142,105,104,99,97,93,111,93,90,90,90,105,106,101,112,104,79,99,99,81,76,99,87,87,89,90,89,74,94,93,93,91,96,88,84,87,87,87,77,97,97,98,100,108,106,106,95,102,99,85,98,98,108,107,98,102,108,105,107,108,75,108,106,106,110,114,117,121,115,117,118,122,120,119,117,120,127,118,120,122,121,130,126,128,134,127,130,127,122,123,121,124,123,120,123,120,123,120,94,118,120,120,122,130,124,117,115,105,99,98,97,99,95,95,103,102,96,95,110,125,122,126,124,131,138,138,122,124,136,129,120,108,138,135,148,177,169,184,188,193,189,161,176,160,185,196,187,188,189,187,193,190,190,195,192,196,192,195,195,193,190,196,189,193,177,193,193,192,195,198,194,196,193,185,172,191,181,191,192,191,196,
27,73,9,3,3,104,56,112,11,79,86,87,30,10,8,8,3,24,41,62,52,55,40,18,56,30,55,68,34,34,15,3,8,16,72,22,28,56,66,38,31,85,96,143,128,138,134,138,136,146,121,172,143,136,136,149,141,144,138,109,156,156,156,160,156,163,159,158,161,164,156,151,146,145,146,137,141,139,148,147,155,131,115,114,125,157,143,125,136,141,145,152,169,182,184,198,201,201,202,201,201,202,211,196,208,202,205,212,207,205,210,210,209,207,208,208,209,209,210,206,207,209,210,210,207,205,209,209,210,207,208,208,206,211,209,210,207,208,213,207,212,214,213,211,211,213,216,212,211,211,208,208,211,209,211,210,210,211,211,210,208,202,214,210,210,210,209,210,211,206,211,209,211,208,210,212,209,208,208,206,204,202,189,197,201,159,202,167,205,170,197,173,194,197,202,201,205,203,202,199,199,198,200,200,203,201,201,199,203,201,201,202,200,200,198,201,202,203,196,194,194,193,192,193,192,194,192,194,195,197,197,191,191,190,196,200,194,199,196,185,192,192,193,188,191,192,192,199,198,194,174,183,190,192,189,187,
153,33,8,1,31,121,170,153,57,21,87,74,70,69,97,131,55,8,7,28,52,16,55,89,12,21,17,29,22,19,23,40,3,36,42,65,132,36,107,14,97,144,181,169,173,204,204,202,206,204,203,202,202,197,201,201,205,201,205,202,203,203,199,202,198,202,201,164,173,196,196,197,198,205,200,196,204,202,206,182,204,204,206,203,202,191,186,193,209,210,205,203,207,205,206,205,208,206,209,212,209,207,211,208,204,201,207,202,205,203,207,208,208,206,206,206,205,207,207,203,205,203,205,205,203,204,201,202,199,202,202,198,203,200,201,202,203,202,202,205,203,205,204,204,206,206,202,200,203,202,202,204,206,208,201,207,206,207,205,204,204,204,203,204,205,207,207,203,204,206,206,205,203,204,204,204,203,204,203,201,203,201,199,200,198,197,199,198,193,190,201,200,201,202,206,199,203,199,200,203,200,201,200,201,199,201,199,200,201,201,200,202,202,200,201,199,198,197,198,197,193,196,196,198,199,196,197,196,195,194,197,192,194,197,196,196,194,197,192,191,195,194,198,199,198,198,195,195,196,196,191,190,191,192,191,193,
92,56,20,1,10,131,141,76,52,5,33,68,28,7,34,103,68,164,76,59,50,31,37,29,38,25,8,12,11,13,43,41,89,48,36,39,45,34,35,13,16,117,138,170,163,188,190,193,190,196,191,190,193,195,192,190,192,191,192,190,194,190,192,195,190,188,188,174,186,196,185,194,193,192,194,197,193,189,80,179,194,193,118,194,197,199,188,202,200,201,191,203,200,200,199,201,202,202,200,201,199,202,201,201,199,199,200,201,203,201,204,201,201,203,203,202,202,201,204,204,202,199,204,199,202,204,202,199,202,201,202,202,201,203,202,201,201,205,203,202,201,202,203,201,204,205,203,205,203,203,204,205,202,205,202,204,207,206,207,206,204,204,200,200,204,205,206,205,204,203,203,204,204,204,204,204,206,205,203,203,202,202,203,201,200,199,200,200,203,200,196,199,199,201,200,202,202,201,199,198,198,201,199,198,198,197,198,197,198,196,195,197,196,198,196,196,197,196,194,196,197,196,195,194,199,197,197,197,196,195,196,197,193,197,194,195,191,193,201,199,197,197,196,194,197,197,197,196,197,194,194,194,192,191,190,189,
16,34,32,5,1,2,16,8,28,9,3,19,18,65,82,115,63,104,17,174,71,45,26,13,13,8,17,16,20,23,16,30,77,22,63,18,8,15,2,11,33,173,97,103,137,190,192,185,192,186,192,190,192,195,196,195,197,197,193,194,196,201,198,199,193,197,200,195,196,194,193,191,190,192,197,191,181,161,181,182,191,183,187,180,177,178,201,196,201,204,203,204,202,203,202,202,201,203,200,204,204,203,206,203,204,202,203,205,201,205,204,203,195,200,204,204,201,203,203,204,203,206,206,202,204,203,203,200,200,203,203,204,204,202,202,203,200,202,201,206,205,206,204,205,206,204,205,204,203,205,208,204,202,203,205,205,203,206,205,202,203,205,202,204,203,203,206,203,204,202,200,204,204,201,201,201,201,198,199,202,203,201,203,202,202,203,202,201,201,196,201,203,202,202,198,194,195,202,204,204,203,201,200,199,199,202,203,203,201,204,200,202,204,202,203,199,203,201,203,202,199,202,201,199,200,203,203,201,202,200,201,201,202,201,201,202,201,203,202,197,199,200,202,201,202,201,201,200,202,201,201,201,200,198,197,198,
6,3,10,2,7,20,5,5,5,8,9,5,9,28,48,63,61,76,39,83,40,51,5,8,7,6,23,48,20,46,65,123,84,36,70,27,21,8,18,8,38,24,22,62,146,192,195,194,193,192,197,194,195,194,197,195,196,197,197,199,192,193,197,195,199,197,199,197,199,190,192,190,196,189,181,188,153,150,153,180,169,165,184,174,164,129,203,203,201,206,204,204,203,206,205,204,205,202,206,203,204,206,206,203,201,204,205,205,204,203,204,201,203,201,207,207,202,203,203,202,203,200,201,202,199,204,198,201,206,201,202,202,200,204,204,202,204,197,205,203,204,202,204,201,206,204,205,204,206,203,204,206,205,203,201,202,203,202,206,208,204,202,204,200,201,206,201,205,201,203,205,202,205,203,203,206,204,205,206,204,203,204,198,205,201,204,202,201,203,201,201,202,200,198,199,201,203,203,202,198,201,203,200,201,202,203,200,202,200,199,199,200,202,201,203,200,203,199,197,202,202,202,200,201,202,202,200,202,199,198,202,200,203,202,200,202,202,202,202,201,198,201,199,202,202,199,196,201,199,200,199,199,199,200,199,195,
3,4,26,4,24,5,4,1,5,12,5,15,6,24,39,26,24,126,138,8,44,64,37,7,9,7,25,18,62,24,109,142,97,82,110,55,26,100,141,23,56,189,187,115,198,194,195,197,195,193,191,192,197,193,196,195,195,196,195,192,194,194,193,195,197,194,197,199,197,197,197,191,192,195,204,194,156,159,173,167,164,166,184,187,189,195,205,200,197,201,197,200,200,197,198,198,200,199,200,201,197,202,204,202,204,195,204,201,206,202,200,201,201,197,202,203,200,203,202,201,199,197,198,202,201,203,200,201,200,199,201,202,204,205,202,203,205,204,205,204,208,204,205,203,205,205,207,204,202,205,200,207,205,203,201,205,203,204,206,205,205,207,201,204,202,202,201,203,203,201,200,199,203,202,199,193,204,201,205,202,198,200,201,203,200,201,202,201,203,202,202,201,202,202,202,202,203,204,204,204,201,203,200,202,202,201,202,200,203,203,200,203,203,196,201,198,200,198,202,201,197,198,199,187,202,200,201,199,200,198,193,204,202,204,197,199,198,195,197,201,193,199,198,198,196,197,195,195,197,197,197,199,200,200,196,194,
3,1,12,3,6,2,2,5,4,5,2,7,7,3,116,32,32,68,110,86,4,42,9,19,13,8,7,10,17,102,91,142,195,103,177,37,54,27,191,140,150,76,147,136,188,193,189,192,192,195,196,196,195,195,195,193,193,195,194,195,193,194,196,194,195,196,197,196,193,195,194,194,195,194,194,202,203,206,203,198,192,196,197,198,200,198,200,199,198,198,199,198,197,198,201,199,200,200,202,199,199,199,202,197,199,201,201,201,201,200,200,202,199,199,201,201,200,200,199,201,201,202,198,197,200,203,200,201,198,201,198,199,200,197,199,199,201,201,201,200,201,200,202,200,200,200,202,199,200,199,199,199,202,202,198,202,201,199,201,203,201,200,198,201,200,199,198,198,195,199,196,199,200,191,199,200,197,201,199,200,201,199,201,200,199,201,200,199,198,199,200,201,200,200,199,198,199,199,194,196,198,197,198,198,198,198,199,195,199,196,198,197,199,199,197,195,197,201,197,195,194,193,193,195,187,189,189,192,193,194,193,193,194,193,192,193,192,192,192,187,195,193,193,194,193,192,193,191,191,191,191,190,191,192,191,192,
1,2,1,1,3,3,2,4,5,5,3,9,8,10,5,4,94,102,163,57,76,3,14,8,5,11,11,10,36,124,102,173,196,143,112,86,96,67,160,189,164,186,127,185,190,188,189,190,191,192,185,189,190,190,192,192,190,191,192,192,191,191,193,191,192,192,192,194,192,190,192,194,191,193,189,191,190,191,186,194,194,196,196,192,199,195,198,197,196,195,196,194,195,193,193,193,194,193,194,195,195,196,195,195,196,196,196,197,196,195,197,196,197,197,196,196,194,195,192,197,195,193,196,194,195,197,193,198,192,193,196,194,192,196,193,195,195,196,198,195,197,193,197,196,197,198,193,198,192,196,196,197,197,196,194,196,193,198,197,195,198,190,195,191,191,194,192,194,195,194,197,197,195,194,193,193,193,193,192,193,196,194,195,195,195,197,194,195,192,194,193,195,194,194,193,192,191,189,192,190,192,193,195,191,191,192,192,190,189,193,186,189,189,187,189,187,187,190,187,187,188,188,188,187,185,187,189,188,188,187,187,183,185,185,183,185,184,183,185,185,185,184,180,182,184,186,184,184,184,186,185,184,183,183,186,184,
4,2,1,2,3,1,4,3,4,5,2,2,22,45,17,10,110,6,73,32,69,15,6,7,9,8,13,25,28,89,156,172,188,168,127,32,121,76,99,175,187,184,179,182,186,184,185,183,184,185,184,186,184,183,184,184,186,186,185,185,184,185,186,186,185,185,186,185,185,182,187,186,184,185,186,184,187,189,188,189,189,188,190,190,188,190,192,186,190,190,188,189,191,188,187,191,190,189,190,191,191,189,193,190,190,193,190,191,189,190,191,188,190,187,192,189,187,192,191,189,193,189,190,191,193,192,192,190,190,187,189,190,190,187,190,188,186,189,191,191,189,187,184,184,191,190,190,191,190,193,191,190,192,188,189,190,193,188,189,188,184,185,188,188,185,186,187,188,186,189,190,188,190,191,188,190,189,192,190,191,188,185,184,185,184,187,185,186,188,187,187,187,187,188,186,188,187,188,187,184,186,188,185,173,176,174,175,181,185,185,185,184,185,185,183,182,182,184,184,185,183,186,186,184,187,183,186,183,185,183,184,180,183,182,179,180,180,181,178,177,179,177,178,176,180,180,179,179,177,178,181,180,180,179,178,182,
0,5,1,1,2,2,7,7,2,15,11,7,30,25,10,2,19,36,19,4,17,6,6,10,12,63,22,27,57,66,147,174,179,177,86,58,70,132,75,182,180,185,180,180,182,178,180,182,179,180,178,181,183,181,180,180,182,180,181,180,178,180,181,181,184,182,183,187,182,183,184,185,184,184,184,184,182,183,182,182,185,186,185,187,186,190,185,186,186,185,185,187,187,183,185,187,189,186,186,188,185,185,186,189,188,186,189,186,184,185,190,186,186,186,186,188,187,188,188,187,183,183,187,188,187,189,187,188,189,189,188,189,188,188,190,188,190,193,189,188,189,185,187,186,189,188,186,188,187,189,185,189,186,187,185,186,184,183,187,186,185,186,185,185,187,187,187,184,189,184,183,184,191,190,189,188,191,194,192,196,194,196,195,203,199,179,182,183,180,184,182,186,182,179,179,177,181,196,196,197,198,198,194,192,197,194,197,198,199,200,193,181,185,182,179,179,181,183,181,180,183,200,201,202,202,202,204,205,205,204,204,207,204,205,204,173,178,178,176,180,179,178,181,181,181,183,200,199,199,199,196,200,199,201,200,202,
1,7,8,4,2,3,2,2,1,1,5,9,2,89,30,8,13,4,4,6,8,4,4,6,6,11,34,29,45,77,96,137,167,181,112,151,141,127,115,176,179,179,182,181,179,178,176,175,180,181,177,180,177,177,178,181,183,195,198,200,200,201,202,200,202,204,203,203,203,186,184,180,178,183,183,180,183,181,179,183,181,208,206,207,204,208,207,207,204,205,186,182,183,184,178,188,187,184,187,184,182,188,208,208,209,211,209,208,209,211,211,208,213,188,186,189,185,187,186,185,184,181,186,184,203,209,215,215,211,212,209,210,212,211,212,201,211,186,187,188,189,184,186,188,188,187,187,188,185,192,190,192,187,188,188,189,189,186,189,190,189,185,187,181,184,183,187,186,185,184,178,183,182,182,186,182,179,179,183,183,181,182,179,179,181,177,181,178,179,182,170,177,178,181,180,181,179,177,174,175,173,170,168,167,173,172,170,165,169,169,170,170,167,172,179,173,176,177,176,179,177,173,177,174,175,175,173,169,173,171,171,174,175,175,176,174,177,174,174,177,171,175,177,173,177,173,176,172,173,172,166,173,172,172,168,173,
0,3,2,2,3,1,2,2,3,4,18,30,26,8,2,2,2,29,3,7,3,5,3,6,1,20,16,32,45,41,122,126,155,170,157,119,183,175,160,177,177,173,177,176,170,175,175,182,177,179,173,171,173,170,172,176,176,172,181,172,178,171,177,176,179,180,184,175,180,177,174,176,178,172,176,178,178,180,177,181,176,176,178,179,179,181,177,177,178,183,181,183,180,180,180,184,181,179,180,184,181,176,184,179,179,187,187,179,180,183,181,181,180,182,177,181,183,183,184,182,184,185,181,185,180,184,188,186,187,185,181,179,178,180,183,186,180,184,179,185,180,179,179,180,179,184,183,180,182,181,185,182,182,183,184,181,183,181,186,183,180,181,180,183,182,184,186,179,182,186,186,181,182,181,178,188,180,181,180,184,180,184,180,177,181,179,177,178,180,182,178,176,176,179,179,177,178,178,175,176,174,176,178,173,174,176,171,175,176,172,171,172,176,173,174,174,172,170,173,176,171,177,175,180,172,170,178,173,176,176,175,175,174,173,173,171,171,167,168,176,171,168,170,166,174,171,173,171,169,171,168,167,166,171,169,172,
2,2,3,2,1,1,4,2,4,1,6,8,43,1,8,2,3,6,1,3,1,4,2,3,15,17,10,15,52,59,131,161,150,164,57,160,152,154,180,173,178,175,172,173,173,176,177,171,174,174,177,175,173,173,173,173,176,176,176,176,177,177,177,175,175,177,174,180,179,177,175,174,173,174,173,173,176,177,180,177,173,178,173,182,181,175,178,176,178,186,172,181,176,177,175,181,181,179,181,180,180,185,179,181,177,177,181,179,180,181,181,182,184,180,177,185,182,178,183,183,170,180,184,181,180,183,181,185,184,181,179,181,178,180,181,179,180,181,176,180,178,183,181,179,177,179,177,175,182,178,185,177,179,187,180,180,181,178,180,183,178,182,180,180,180,176,180,179,179,180,178,179,180,178,179,178,175,180,176,177,183,179,180,177,178,177,177,171,174,171,172,173,173,173,175,174,173,176,173,173,173,175,172,173,174,174,174,171,173,172,173,169,171,166,163,169,168,169,172,167,171,167,169,168,166,162,168,167,167,169,159,171,171,160,163,164,168,164,166,163,160,161,164,167,154,164,160,164,161,159,167,160,158,158,158,165,
1,1,1,1,1,1,1,3,0,1,8,1,11,21,5,2,2,1,2,2,2,2,1,2,6,5,7,14,27,46,104,98,150,165,172,172,165,167,163,172,170,173,168,170,171,166,171,168,170,172,169,171,167,166,167,168,170,169,164,171,170,166,169,169,168,177,177,169,174,171,173,172,173,176,175,173,174,180,173,176,177,173,175,177,172,180,173,177,179,179,178,179,181,176,178,176,177,176,181,174,173,178,178,178,182,177,174,180,174,179,183,178,179,181,179,180,176,177,177,179,183,171,180,179,181,179,175,178,178,175,175,169,179,174,181,178,179,180,174,179,181,174,175,177,177,177,173,181,179,183,178,179,179,182,177,174,175,180,180,175,177,181,180,177,175,176,174,174,176,174,175,177,176,176,177,175,177,178,171,176,176,177,176,172,175,176,170,173,174,175,175,172,173,174,172,174,172,174,172,174,169,169,166,168,169,171,169,166,168,169,165,168,165,167,172,166,165,168,169,165,166,167,162,167,165,167,162,162,164,161,162,162,162,164,166,162,159,164,164,165,163,160,164,160,159,163,167,161,165,157,166,163,157,161,158,159,
0,0,1,1,1,1,1,1,0,1,2,7,15,0,4,2,2,1,2,0,1,1,1,0,7,4,5,8,44,76,88,136,151,68,173,171,172,167,167,163,169,168,172,167,167,167,165,168,169,168,165,166,166,168,164,172,168,169,171,164,169,167,168,167,168,170,172,169,167,171,164,172,171,168,173,168,171,171,168,172,169,173,167,172,170,175,173,167,172,174,169,173,171,169,171,174,175,175,172,176,174,174,173,174,171,167,176,174,173,174,176,177,176,178,176,174,172,176,178,174,179,171,173,174,175,175,178,177,170,178,173,170,174,173,176,169,174,177,176,180,176,173,177,177,174,175,175,175,180,179,179,175,176,179,179,178,179,177,177,178,182,180,175,177,177,183,175,173,178,175,177,176,173,174,176,173,173,173,176,170,181,174,172,174,175,170,175,173,164,173,172,165,175,173,170,173,169,168,175,169,172,169,170,170,173,169,170,165,169,166,167,166,165,165,165,166,168,166,167,160,161,161,164,164,166,169,165,167,164,166,164,166,163,162,161,162,165,162,161,160,159,158,159,157,153,152,156,158,155,155,162,158,158,155,154,155,
0,0,2,1,1,0,2,1,2,1,1,12,3,10,3,3,4,0,1,0,0,0,1,2,2,2,5,10,8,38,49,131,143,167,174,168,169,167,167,169,169,167,167,167,165,166,169,167,164,169,164,167,171,167,166,170,174,168,172,170,167,169,174,175,176,172,175,170,168,170,168,170,171,173,172,170,170,168,170,170,167,167,168,168,173,170,168,172,171,168,170,168,170,166,166,171,170,172,174,168,171,168,171,174,171,177,174,176,176,172,173,174,177,173,177,175,172,172,172,175,173,167,172,174,177,168,167,165,171,172,168,168,171,171,172,172,172,172,175,167,174,171,167,173,169,174,175,174,176,171,167,176,175,175,180,177,175,175,173,171,173,170,174,172,169,170,171,170,169,174,172,169,167,173,172,171,170,175,171,171,176,160,170,172,171,167,171,171,174,173,166,171,167,169,161,167,168,168,170,168,162,172,171,170,172,168,163,167,169,166,169,167,170,164,167,167,167,170,168,165,161,167,165,164,164,157,159,167,156,168,164,163,163,157,163,164,163,161,164,162,164,160,157,160,164,150,158,155,155,151,161,158,157,158,158,156,
1,1,0,2,1,1,2,1,4,1,10,3,11,3,0,0,1,0,0,0,0,2,1,1,3,1,2,5,20,63,156,107,56,166,170,175,168,169,167,167,167,168,167,165,164,161,167,164,167,167,157,159,165,162,169,164,168,169,170,166,169,166,171,168,168,169,166,168,164,170,165,167,164,162,169,169,170,166,165,168,168,164,170,166,172,171,169,167,171,161,168,174,170,171,170,166,169,171,172,170,171,172,169,172,167,170,170,168,169,172,174,175,170,171,170,170,168,166,169,169,170,174,171,171,170,173,168,168,167,170,167,174,176,173,171,170,169,169,167,170,170,173,169,173,173,172,173,171,171,169,175,172,174,168,171,171,169,167,176,169,172,170,176,172,169,170,159,165,168,172,171,169,171,177,170,174,172,172,172,172,168,173,169,172,172,171,171,171,175,174,175,171,171,175,171,176,174,168,179,172,169,173,177,175,171,166,163,167,172,173,172,170,169,171,167,170,174,172,166,170,166,169,171,174,156,173,166,168,164,171,163,162,166,162,164,167,164,163,172,164,165,162,161,165,157,160,147,161,163,172,160,162,161,159,166,161,
2,1,2,1,1,2,2,1,1,5,3,1,5,1,0,0,1,1,0,0,2,0,1,2,2,3,8,29,107,172,162,8,169,173,168,170,166,168,176,169,169,169,167,166,163,167,168,167,160,160,176,164,165,164,168,165,167,170,163,167,167,169,171,173,168,170,166,168,169,168,172,169,167,163,166,171,171,164,167,166,169,169,171,171,170,171,171,167,169,170,167,172,170,167,167,167,171,173,171,168,169,162,161,166,169,168,172,170,168,168,168,168,172,170,167,173,171,176,173,174,170,170,175,168,170,169,172,166,172,176,171,171,169,167,170,179,176,177,167,172,174,170,169,175,170,170,168,169,166,174,172,172,170,169,171,174,174,173,178,172,174,173,174,179,173,176,176,170,174,178,172,182,179,178,180,179,172,183,174,177,178,178,175,176,179,177,174,181,176,180,183,179,175,176,176,181,173,176,175,171,178,180,175,167,170,172,174,172,180,174,176,176,177,179,174,177,177,171,178,177,174,169,176,173,174,172,174,176,171,176,168,174,172,173,174,172,168,172,176,176,178,173,175,171,167,162,170,172,169,170,167,168,170,165,162,168,
5,5,1,1,1,1,3,4,1,1,1,0,0,0,1,1,0,0,0,1,0,1,1,3,8,6,24,69,143,80,42,167,173,171,166,170,170,169,170,170,167,170,171,167,169,167,169,167,168,171,172,173,173,171,172,172,172,171,175,171,173,169,173,168,172,173,168,170,173,172,176,173,172,173,173,172,176,170,179,179,175,175,170,176,173,172,178,168,171,171,175,174,171,175,175,179,177,181,177,173,173,173,171,179,178,177,178,178,180,180,178,178,177,176,179,176,183,179,182,179,179,186,181,179,182,181,176,177,176,176,174,176,175,173,176,174,179,177,178,175,176,178,179,178,177,180,177,177,182,177,179,184,178,182,176,180,178,173,175,179,175,175,182,179,179,173,175,177,177,180,179,178,175,176,179,174,178,177,176,176,185,183,183,174,176,178,176,176,176,183,176,176,177,176,174,176,177,174,170,173,171,174,177,177,175,165,170,170,173,175,173,175,178,175,173,173,171,177,179,183,173,174,175,172,173,169,172,171,175,173,170,174,168,166,167,169,178,174,175,170,172,173,172,171,172,173,173,171,168,167,167,155,169,168,169,166,
2,1,2,0,0,0,0,3,1,1,1,0,1,1,1,0,0,0,0,0,1,1,3,5,5,24,89,100,16,156,170,176,172,169,170,172,168,173,170,166,171,167,167,168,170,169,173,168,172,170,165,166,167,169,170,166,168,168,170,174,169,174,168,173,174,167,169,173,175,169,175,172,176,169,173,173,177,173,176,180,179,177,173,177,173,176,176,176,172,183,180,173,179,168,176,179,178,176,174,178,179,179,178,178,180,180,180,180,176,179,177,180,177,176,175,175,180,175,175,177,181,175,180,177,180,179,178,180,183,176,181,178,175,177,175,178,179,175,186,174,177,180,179,177,178,185,178,174,179,184,179,183,187,181,184,178,179,180,183,179,184,180,182,178,183,173,181,178,181,177,183,176,176,177,176,178,177,176,175,176,178,184,187,178,182,177,173,175,177,178,175,175,181,178,179,180,176,175,175,172,180,175,174,178,177,174,175,175,177,175,180,176,182,175,168,175,175,174,175,175,193,175,174,176,181,177,175,178,172,173,168,177,177,166,170,173,169,175,166,172,169,169,175,167,170,168,172,171,174,171,167,171,169,168,169,166,
20,3,5,1,1,0,0,0,0,0,0,1,1,0,0,0,0,0,1,1,1,1,4,18,6,87,25,75,135,162,137,174,174,173,173,166,174,161,169,168,174,173,169,172,173,173,169,164,174,167,169,170,176,171,164,170,174,170,169,174,176,170,173,172,168,172,168,176,173,172,171,174,172,179,173,173,174,166,173,175,177,174,177,176,169,172,168,170,171,173,176,176,174,178,174,178,174,170,173,169,172,176,178,177,177,178,171,170,178,174,178,171,176,176,180,176,180,182,175,177,175,185,180,180,177,179,175,184,182,174,178,176,175,178,183,180,174,182,184,171,178,181,181,176,177,181,178,178,180,179,179,184,184,181,186,184,180,182,178,173,180,174,178,180,177,176,176,173,177,181,180,176,175,175,176,173,171,174,178,172,174,173,175,174,174,182,180,176,174,176,171,184,179,177,175,174,176,182,169,174,174,172,176,173,174,172,175,176,174,175,178,172,173,173,168,176,175,176,178,175,176,175,168,174,171,171,175,172,176,173,177,169,173,179,169,168,173,170,168,169,169,168,170,169,168,170,164,170,170,167,168,171,167,165,163,166,
17,4,2,0,2,2,13,0,0,0,0,0,0,0,0,0,0,0,1,1,3,2,50,18,23,4,48,142,115,158,169,167,169,173,167,166,166,169,165,166,167,164,167,171,171,170,167,167,168,168,169,163,165,165,162,163,166,164,167,168,168,171,167,163,173,167,166,168,169,170,171,170,172,176,172,172,168,171,176,171,173,176,170,174,172,177,186,176,174,175,170,181,176,175,171,180,174,173,173,174,175,172,186,177,178,180,176,173,171,177,179,179,178,181,176,180,177,175,176,181,174,179,173,182,180,180,174,180,180,178,177,175,184,180,181,181,178,181,176,176,180,175,179,179,176,175,179,176,177,178,180,181,178,178,181,184,179,180,180,185,188,182,180,181,181,180,177,184,180,179,183,176,179,177,180,182,177,176,178,179,177,181,176,176,179,176,178,177,177,178,177,175,181,180,181,173,173,177,179,176,174,173,175,175,175,176,176,177,176,174,175,182,174,178,179,176,176,172,176,175,176,170,176,178,176,175,175,181,178,176,175,173,174,174,173,174,171,175,171,179,175,174,170,168,176,160,176,171,173,179,168,171,173,169,173,167,
9,17,1,0,6,2,10,3,1,1,1,1,1,1,1,1,1,0,1,1,1,1,2,2,19,38,104,120,155,120,149,160,172,173,171,171,172,170,168,168,170,175,173,174,169,168,172,169,172,171,169,172,169,169,167,176,175,173,172,172,174,174,171,178,173,178,179,171,172,171,167,176,172,172,177,174,178,170,172,178,180,176,185,177,174,170,180,177,178,181,173,176,176,173,177,174,177,172,178,179,183,180,184,178,175,178,176,181,178,179,181,180,182,180,182,183,179,182,177,179,178,186,178,178,183,184,178,176,184,179,181,180,180,182,181,183,176,180,182,183,183,183,179,179,181,178,185,177,182,179,181,176,180,185,181,179,178,187,179,184,181,175,184,187,188,178,176,181,175,187,179,185,184,184,178,181,183,171,176,180,187,180,179,179,177,171,173,180,178,178,180,180,174,175,181,179,179,179,177,178,180,177,173,180,179,178,175,178,178,176,181,179,180,179,175,180,180,178,175,178,177,175,175,180,176,180,178,178,175,181,175,173,175,171,174,178,177,177,172,178,172,175,175,178,175,176,176,175,172,177,172,170,168,171,170,172,
27,5,5,2,3,3,0,3,1,7,0,7,2,3,0,2,4,0,2,1,0,7,8,136,105,43,147,127,107,101,146,176,179,173,174,174,176,173,174,173,171,169,178,173,176,177,173,172,172,171,170,177,154,119,175,166,180,169,178,179,172,171,179,169,171,178,172,179,177,174,182,178,174,185,178,177,176,180,180,181,180,183,179,182,175,168,182,180,181,179,185,182,181,181,186,182,179,183,183,181,182,180,181,180,181,185,174,186,183,178,179,183,183,179,181,179,183,181,177,184,184,180,175,182,178,180,178,186,179,185,182,182,174,181,180,182,190,186,178,182,181,182,185,192,183,184,184,181,184,182,177,181,183,184,177,167,175,183,181,182,184,182,189,185,185,183,187,181,184,188,186,185,183,180,187,182,175,175,180,188,184,183,174,180,180,185,158,174,186,186,180,187,181,182,177,181,182,179,180,181,177,179,177,177,183,179,177,179,189,179,179,180,181,179,182,179,176,177,178,182,176,174,174,174,180,179,183,175,180,179,180,175,176,187,181,177,175,178,179,173,175,176,179,175,180,178,177,180,177,177,180,176,177,174,176,176,
3,3,0,2,7,4,2,2,0,17,5,24,20,4,3,12,2,6,2,1,2,13,100,174,156,108,18,168,183,179,180,175,171,181,174,176,178,180,182,174,176,177,179,175,176,162,162,168,170,170,130,135,131,112,86,169,178,177,174,179,183,181,177,181,183,180,180,178,180,188,186,182,181,176,184,178,183,183,183,184,182,179,183,185,184,180,179,182,178,181,185,184,182,184,180,181,179,183,185,181,178,191,180,188,183,186,185,179,180,184,189,184,182,182,186,190,184,184,185,184,187,187,178,182,189,183,182,182,184,185,184,180,184,186,185,181,184,179,186,181,183,186,184,184,184,187,189,187,186,188,187,184,184,188,189,182,188,192,191,185,182,184,181,189,186,182,186,182,189,182,187,184,181,183,186,185,190,187,188,186,185,178,187,179,185,187,181,185,185,181,183,185,181,179,182,182,181,182,182,183,182,182,182,181,179,202,205,204,202,202,204,202,202,203,204,202,202,202,201,203,202,203,200,201,204,201,203,201,200,200,197,199,201,199,201,203,199,196,201,192,199,195,197,196,197,197,194,194,179,181,178,180,178,181,177,173,
1,1,2,1,1,3,7,9,2,5,25,27,6,8,1,4,7,4,4,42,48,16,39,15,25,109,129,119,151,149,183,175,182,181,178,178,178,181,176,183,180,186,182,189,186,185,186,184,191,111,98,78,74,111,55,188,193,199,199,198,202,199,198,201,197,204,204,202,203,201,203,202,201,201,184,176,183,183,181,181,185,182,182,181,183,182,180,183,181,187,180,180,188,185,183,184,190,190,188,189,186,185,186,189,189,182,183,188,184,186,190,187,189,185,189,181,188,205,210,206,203,210,209,208,207,207,206,207,204,204,201,196,192,189,192,192,195,189,194,196,193,196,193,197,196,192,197,195,194,194,193,194,194,193,190,190,177,188,184,192,188,193,183,189,186,183,183,187,188,187,188,187,188,189,186,184,187,184,187,184,180,186,189,191,186,193,184,189,193,183,186,184,183,179,185,185,183,184,188,187,181,187,187,187,187,179,179,180,179,178,182,177,182,186,177,179,178,182,185,187,180,178,176,176,178,177,180,178,178,181,177,181,179,178,177,182,180,178,179,178,181,177,180,177,176,179,180,180,179,180,182,177,175,172,172,170,
4,12,1,1,1,5,12,54,16,3,3,2,1,3,6,12,25,6,20,25,21,7,75,110,53,60,103,124,151,184,180,177,179,176,181,176,176,175,188,191,190,182,190,189,190,187,189,187,181,124,38,53,95,115,109,111,179,177,184,177,181,181,179,180,184,180,173,184,179,180,179,182,184,178,180,182,183,182,180,185,180,177,177,179,178,183,181,183,185,179,182,188,189,183,182,183,189,181,179,186,183,182,184,185,186,187,185,186,179,184,186,184,183,185,186,185,186,183,185,187,189,190,185,184,190,187,184,181,190,186,182,188,186,183,188,186,190,187,184,189,191,185,187,177,185,183,186,183,186,185,191,189,191,191,187,190,194,192,191,189,191,187,189,188,184,186,178,191,190,188,188,190,185,190,194,192,189,192,191,186,184,189,188,188,187,186,185,182,183,184,183,180,180,183,180,182,180,173,178,180,182,180,179,183,180,179,181,176,179,177,180,176,176,179,179,181,175,179,175,181,182,177,175,175,179,176,175,176,177,178,178,175,177,172,175,175,175,178,174,176,175,173,175,171,168,173,175,166,170,171,170,174,171,172,171,174,
2,6,3,1,1,3,2,4,6,8,19,3,17,13,59,8,65,56,107,55,25,61,19,8,44,120,126,155,147,183,177,176,174,180,181,176,181,172,167,178,176,175,177,175,175,184,176,178,172,138,10,44,110,106,54,117,173,180,174,175,179,176,178,175,174,179,176,173,179,177,176,177,176,178,177,179,181,177,181,181,178,179,182,175,179,180,176,184,173,182,178,183,177,165,187,180,184,183,180,185,180,178,184,182,183,183,184,183,186,184,187,178,182,185,183,182,185,186,180,186,182,185,180,185,188,189,186,180,185,183,191,183,182,182,183,182,181,182,181,181,186,182,182,187,183,181,182,182,182,186,187,184,186,183,183,186,178,181,183,184,182,180,183,187,187,183,185,184,182,185,184,184,182,188,184,184,177,181,197,185,185,184,179,183,182,183,185,179,179,182,180,188,175,186,182,179,178,180,188,184,182,181,186,178,180,179,182,179,173,172,183,177,183,179,177,181,177,179,178,180,176,177,167,174,178,169,175,171,174,178,171,175,173,173,175,177,172,174,174,177,170,175,170,166,170,170,167,169,169,170,167,167,167,168,168,168,
0,2,1,2,0,1,6,58,32,28,11,4,6,43,25,30,23,42,84,95,67,35,19,33,31,41,120,178,180,178,177,171,179,177,175,179,177,177,167,176,174,175,175,177,182,177,174,172,172,92,19,57,28,37,86,176,178,171,177,182,178,183,175,172,176,176,174,181,175,180,179,180,180,179,181,180,179,183,178,182,178,182,182,178,183,181,180,183,175,175,177,184,179,176,181,178,184,184,186,182,182,187,184,181,181,179,180,182,187,188,183,181,183,183,184,186,180,184,188,185,183,179,185,179,180,184,181,178,188,185,181,180,177,178,181,182,171,171,186,185,182,181,178,182,183,181,186,184,182,175,172,184,179,186,173,185,184,189,183,185,178,184,181,179,183,183,181,180,184,183,180,180,186,185,181,180,183,181,178,179,183,184,182,180,183,176,180,182,180,176,181,180,177,178,176,177,174,185,178,180,180,174,177,176,179,171,174,176,177,171,171,172,172,174,174,180,174,172,169,176,172,170,165,171,167,166,171,167,169,166,164,171,175,169,174,172,169,165,168,169,169,167,168,161,170,159,156,167,164,159,163,165,166,163,166,161,
1,0,0,0,3,2,6,6,5,1,4,3,41,88,81,75,87,93,50,81,77,55,21,7,52,44,91,155,147,182,168,153,172,173,179,174,174,176,182,175,173,184,171,173,169,174,177,170,108,87,10,28,27,6,49,176,171,172,175,170,171,172,174,174,181,173,181,179,173,165,174,174,169,170,174,174,177,180,175,172,176,175,174,174,179,178,171,174,178,186,185,178,180,180,183,186,173,177,175,179,181,177,183,181,184,183,180,176,178,186,181,172,177,174,181,179,176,181,175,178,181,172,180,184,177,175,180,177,176,178,178,176,182,181,180,176,180,185,177,177,177,177,177,177,180,183,184,183,183,174,184,182,183,178,176,183,177,177,172,180,182,171,177,177,175,169,174,178,176,176,176,173,172,169,178,182,178,179,173,174,173,179,171,168,177,171,181,175,171,176,170,175,176,174,177,179,170,170,178,169,173,174,176,176,168,182,170,176,176,173,170,165,168,169,169,168,170,170,169,169,174,171,163,169,173,170,164,169,166,163,165,162,168,177,161,167,165,164,169,160,169,166,166,158,168,163,157,160,164,163,166,163,163,164,158,165,
0,2,0,0,2,2,3,13,4,0,3,3,55,26,48,115,144,8,14,37,63,28,7,78,18,114,104,76,43,68,45,87,152,155,145,168,168,167,165,157,166,175,173,174,170,165,172,176,167,27,15,5,42,4,23,167,172,168,171,169,177,173,170,165,177,174,163,170,174,176,172,177,167,166,180,170,169,176,181,177,169,169,188,172,183,178,181,174,179,165,165,180,158,175,174,181,172,164,174,169,174,175,176,179,173,174,182,179,172,182,180,180,173,176,178,176,171,177,173,177,177,181,176,181,177,179,181,180,174,179,173,180,179,179,180,170,181,179,179,176,175,184,184,172,177,176,176,163,179,181,178,178,177,174,173,171,170,186,174,176,170,179,167,175,169,181,182,169,174,169,169,168,176,171,181,183,181,181,180,176,179,172,179,174,176,170,176,177,174,176,171,176,167,171,177,172,159,174,168,179,172,173,166,168,172,167,172,173,172,174,168,165,158,165,168,166,170,168,168,173,165,167,165,170,169,173,161,172,168,168,167,157,169,162,169,168,167,166,158,159,160,159,166,164,156,169,156,162,165,172,167,163,162,161,159,162,
1,2,2,1,2,3,2,1,4,0,2,9,19,24,21,34,54,72,14,5,33,4,5,68,27,83,38,31,50,42,54,116,87,143,163,164,168,173,116,124,152,167,169,166,170,177,169,149,135,22,10,3,7,9,131,170,138,175,169,172,181,177,178,174,175,169,173,170,172,175,176,170,170,180,172,169,182,180,175,178,181,175,175,177,176,170,180,174,173,175,177,178,176,175,187,176,176,175,180,174,173,174,176,174,172,178,171,177,179,177,177,171,180,169,174,169,175,177,177,171,177,173,179,175,174,176,177,174,175,172,182,177,175,172,172,177,174,174,178,164,171,176,172,173,171,170,169,168,176,177,174,177,171,170,174,172,177,175,173,175,171,167,172,175,165,174,182,176,180,179,169,172,164,174,176,176,171,176,171,171,177,174,172,170,173,174,179,173,162,176,174,175,169,173,168,175,171,173,177,173,173,171,172,173,167,173,170,178,168,171,170,170,168,172,168,171,170,172,170,162,168,165,172,167,167,162,170,168,171,164,173,161,164,162,169,164,158,165,164,166,165,164,160,168,167,166,160,168,158,163,162,165,162,153,160,162,
1,2,0,2,0,1,0,0,1,1,1,4,6,9,15,21,33,13,6,8,13,8,16,5,8,61,22,18,15,67,95,43,68,127,174,104,112,100,97,104,160,166,167,172,166,165,166,167,132,20,4,4,28,14,168,170,172,178,170,171,173,163,167,169,170,170,174,173,172,168,167,168,172,167,167,175,175,168,169,171,166,171,170,173,174,172,173,175,173,168,171,174,176,166,177,178,176,178,175,175,179,179,173,180,174,172,166,175,180,179,171,173,169,170,178,177,174,164,171,174,171,180,174,173,178,178,171,173,167,173,176,169,174,176,173,175,170,175,174,168,172,171,175,172,176,175,171,174,175,178,175,180,176,179,173,174,175,170,171,174,171,166,175,179,177,172,180,176,174,167,176,172,170,153,168,170,172,175,174,169,172,169,173,176,181,167,172,173,176,179,170,172,171,170,171,172,172,172,169,176,177,172,172,178,169,174,173,169,172,166,164,172,171,170,166,168,166,172,174,168,167,170,169,169,166,163,169,167,166,164,166,165,163,162,161,166,167,163,159,165,167,164,166,161,162,161,165,158,157,162,164,160,159,153,160,158,
1,2,2,0,3,1,2,1,1,0,1,8,7,9,10,7,19,23,11,8,10,9,4,8,9,5,14,10,15,29,22,24,62,148,37,62,104,15,45,124,144,164,168,169,164,168,169,167,96,11,12,2,24,27,90,152,149,174,168,169,172,176,164,170,170,174,176,173,169,176,173,171,168,172,172,171,160,170,170,172,167,168,168,163,166,175,164,166,165,172,170,171,172,172,173,177,175,174,173,178,174,177,175,178,170,172,173,175,174,178,176,172,174,175,172,174,178,174,172,174,177,179,174,177,176,177,174,176,174,176,176,175,175,177,176,167,170,175,177,174,173,170,170,172,173,169,172,171,177,174,166,164,175,178,173,171,174,177,172,175,173,162,172,174,167,175,174,174,169,175,173,174,177,171,171,164,159,168,165,173,173,174,169,172,175,182,175,172,171,170,175,172,175,178,172,169,168,169,176,166,171,175,168,170,172,167,170,164,165,169,167,162,164,169,165,171,172,170,169,171,163,169,167,166,168,165,169,167,170,170,169,162,164,156,161,161,163,164,168,163,161,162,164,162,160,163,169,159,164,158,158,159,164,168,160,158,
1,1,2,2,2,2,0,0,1,1,0,2,7,4,8,10,9,15,10,13,20,16,25,4,10,5,8,14,3,21,36,15,42,46,49,85,15,19,26,127,121,153,171,170,167,167,171,172,136,7,42,5,13,110,145,165,171,168,180,172,174,170,172,171,178,178,170,168,171,169,175,176,169,174,170,174,175,168,170,170,174,172,176,169,173,170,169,172,173,165,158,167,165,156,174,171,176,171,175,175,175,181,187,174,176,176,180,174,172,172,175,176,176,171,176,173,173,172,175,178,175,179,177,173,177,173,171,181,179,175,173,183,176,178,172,174,173,177,180,174,171,173,174,175,171,177,175,179,173,177,174,179,171,174,172,172,171,175,167,176,170,173,177,170,165,173,168,171,176,172,172,174,179,176,175,177,176,166,170,176,166,168,171,160,171,174,176,171,172,174,176,167,173,169,167,171,175,170,163,168,167,177,175,171,173,176,172,160,174,165,164,172,173,158,168,167,168,162,168,176,168,168,166,167,158,166,153,164,167,166,168,166,166,159,163,161,156,160,159,165,159,157,158,157,165,160,163,161,164,160,159,165,161,162,159,156,
1,1,1,1,1,2,1,0,2,0,4,2,2,4,5,5,12,16,13,10,9,7,12,12,5,7,11,6,11,19,13,11,21,35,10,36,8,9,30,62,86,131,147,163,157,166,172,169,178,21,17,17,18,101,140,169,169,172,172,172,170,167,171,172,164,173,164,166,169,170,133,171,165,151,170,168,167,165,162,170,172,167,169,167,166,170,166,162,167,171,172,170,166,155,143,143,174,168,177,175,176,174,173,174,172,124,167,176,171,175,176,193,182,173,170,171,174,169,176,177,179,184,178,175,174,177,180,181,175,178,180,168,173,173,177,175,179,173,169,174,175,169,174,175,177,172,179,173,175,170,168,166,173,176,176,177,176,169,147,170,177,176,160,169,179,167,171,177,174,172,167,172,167,172,165,172,169,166,176,163,167,175,159,168,169,181,166,177,176,176,173,170,170,170,167,158,173,179,171,169,166,176,173,169,161,167,168,165,167,169,166,171,167,157,167,169,165,170,163,166,169,163,172,160,166,159,161,165,163,168,159,161,157,167,163,166,168,162,166,168,161,167,164,161,158,163,163,162,163,163,156,167,166,164,164,164,
2,2,2,2,1,0,2,1,8,3,3,3,6,6,5,6,9,9,11,9,5,3,6,3,3,13,14,6,8,12,13,12,83,6,3,7,4,15,6,20,63,75,102,134,90,79,148,157,176,7,7,28,79,80,165,168,166,169,171,171,168,172,168,169,170,172,174,174,173,168,175,172,169,170,179,170,174,173,170,172,171,170,178,166,173,178,172,168,175,169,170,173,169,168,177,172,166,182,175,178,178,180,171,174,176,170,173,176,177,174,173,178,175,162,172,181,175,171,144,175,177,181,188,186,198,187,183,191,184,198,180,171,179,168,174,187,174,179,172,171,174,171,176,175,178,177,164,175,172,174,176,172,175,176,174,174,180,174,173,171,166,174,174,170,173,179,180,173,172,172,176,172,177,171,172,171,168,174,166,170,163,174,162,170,169,160,172,165,171,171,173,174,165,171,177,172,170,170,173,182,180,169,168,169,164,176,169,170,168,168,167,165,167,158,170,164,172,169,169,164,167,166,171,170,169,173,169,165,170,163,163,166,168,171,163,168,172,171,166,167,161,163,169,170,169,166,164,160,168,169,164,166,168,168,170,161,
1,1,3,2,4,6,3,2,0,0,4,6,6,4,3,6,10,9,8,1,5,31,1,14,4,7,13,16,18,15,5,9,31,7,4,1,9,11,15,83,32,136,96,17,52,115,102,167,138,65,4,10,73,170,173,169,171,167,169,168,166,171,167,173,174,171,177,169,172,177,174,173,170,175,164,173,168,170,172,174,177,172,170,176,171,164,161,172,172,179,174,172,179,175,176,174,172,178,180,182,177,173,177,175,172,178,174,171,180,175,175,173,179,170,177,178,174,180,174,177,173,168,177,182,178,195,188,187,188,183,184,173,171,171,172,166,173,184,172,174,180,176,177,165,179,175,175,171,178,185,174,167,176,166,167,177,175,177,171,171,171,174,179,174,175,177,178,180,179,177,175,179,174,168,175,180,172,179,176,169,175,174,174,177,181,184,177,173,177,170,177,174,174,179,179,174,178,175,177,177,185,179,184,183,175,170,178,169,174,173,170,177,176,180,179,164,174,173,164,171,176,165,174,169,171,174,170,177,176,178,176,176,176,168,174,169,167,171,168,167,169,165,176,172,167,172,163,162,166,163,169,162,163,168,170,170,
1,1,1,2,2,9,11,6,8,3,7,6,8,4,17,7,6,6,4,5,45,27,4,3,3,9,28,21,15,4,25,35,9,3,3,5,12,12,16,18,14,45,63,62,9,93,107,53,9,75,5,47,171,174,166,170,169,172,174,175,167,174,170,172,169,176,178,179,172,171,171,178,176,174,166,172,172,174,176,180,181,170,175,174,179,170,170,174,179,170,176,171,178,175,176,179,172,177,172,176,180,184,182,180,176,178,179,181,179,180,176,178,178,174,180,178,171,185,176,182,177,178,182,182,177,178,180,183,181,178,179,179,184,178,187,181,182,177,181,178,179,182,185,185,180,178,184,179,180,175,181,186,185,178,186,183,180,176,172,177,177,184,180,177,178,183,182,179,180,174,187,177,179,182,181,182,178,180,181,181,176,181,181,177,186,180,182,179,178,182,173,174,178,186,182,177,173,175,172,175,183,179,180,181,176,176,180,176,179,170,176,171,172,167,172,169,171,172,181,174,167,175,167,173,175,168,175,170,173,172,175,170,177,164,175,173,176,173,172,166,169,169,166,168,170,171,168,166,168,164,166,168,161,167,170,166,
3,0,1,5,2,1,13,22,12,4,11,2,9,3,6,7,8,8,17,14,7,3,5,2,8,13,32,15,34,15,5,4,2,0,3,5,10,9,9,8,10,5,19,32,39,101,136,116,6,5,25,169,170,174,176,176,172,174,174,177,177,183,175,174,172,179,173,179,173,173,176,176,172,171,176,176,172,176,175,176,174,178,176,174,177,180,169,177,182,178,172,176,176,173,179,182,177,180,175,180,178,184,174,181,180,178,177,179,183,184,184,181,183,185,179,189,178,176,181,176,180,182,182,177,176,180,178,178,180,184,177,180,180,182,175,175,176,179,181,186,180,178,177,183,175,183,179,177,182,172,178,183,179,181,176,177,177,179,186,170,179,175,181,175,180,176,182,172,182,175,176,177,174,163,179,183,175,178,182,188,182,182,178,180,178,177,178,174,179,176,181,183,175,182,179,171,179,179,178,176,175,171,173,174,172,176,178,177,174,175,173,176,175,172,177,173,171,176,175,173,166,175,173,175,174,177,174,165,172,165,175,174,173,171,167,172,167,164,166,173,168,163,166,167,168,167,171,168,165,167,168,167,166,170,167,165

);
constant ROM_Gauss: Array4096 :=(154,154,154,154,154,154,154,154,154,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,156,156,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,154,154,154,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,156,156,156,156,156,156,156,156,156,156,157,157,157,157,156,156,157,157,157,157,157,157,157,157,157,157,157,157,158,158,157,158,158,158,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,157,157,156,155,155,155,155,156,156,157,157,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,160,160,161,161,161,161,161,160,160,160,160,160,161,161,160,160,159,156,152,153,156,158,156,149,142,141,143,141,139,
154,154,154,154,154,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,155,156,156,156,156,155,155,155,155,155,155,155,155,155,155,155,156,156,155,155,155,155,155,155,155,155,155,155,155,155,156,156,156,155,156,156,156,155,155,156,156,156,156,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,158,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,157,157,156,155,156,156,156,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,158,154,154,157,160,160,156,149,146,146,145,143,
155,155,155,155,155,155,155,155,155,155,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,155,155,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,155,155,155,155,155,155,156,156,156,156,156,156,156,156,156,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,158,157,157,157,157,157,157,157,157,157,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,161,160,161,161,161,161,161,161,161,161,161,162,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,157,156,158,163,166,164,158,152,151,150,150,
155,155,155,155,156,156,156,156,156,156,156,157,157,157,157,157,156,156,157,157,157,157,157,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,156,156,156,156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,159,159,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,158,158,158,157,157,158,158,158,158,158,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,160,157,154,156,159,160,162,166,167,161,152,148,150,150,149,
156,156,156,156,156,156,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,159,159,159,158,158,158,158,158,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,162,162,161,161,161,162,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,164,163,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,161,157,147,139,145,158,164,165,165,161,147,136,137,144,146,145,
156,156,156,156,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,157,157,157,158,158,158,157,157,157,158,158,158,158,158,157,157,158,158,158,158,158,158,158,158,158,158,157,157,157,157,157,157,158,158,158,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,163,162,163,163,163,163,163,163,163,163,163,163,163,163,162,161,161,160,153,139,131,141,158,165,164,163,155,138,127,134,143,147,148,
157,157,157,157,157,157,157,157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,163,163,163,163,163,163,163,163,163,163,164,164,163,163,163,163,163,163,163,163,164,164,164,164,164,163,162,160,158,156,150,140,138,149,161,164,163,162,155,140,132,136,144,149,152,
157,157,158,158,158,158,158,158,158,158,158,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,158,158,158,159,159,159,159,158,158,159,159,159,159,159,159,159,159,159,159,158,158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,161,161,161,162,162,162,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,163,163,164,164,164,164,164,164,164,164,164,164,163,163,164,164,164,164,164,164,164,165,164,164,164,164,162,160,156,153,149,146,150,159,164,165,163,163,159,148,137,132,133,139,143,
158,158,158,158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,161,161,161,161,161,161,161,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,164,164,164,164,163,163,164,165,165,164,165,165,165,165,165,164,164,164,165,164,164,164,164,165,164,163,163,163,164,165,164,162,158,154,153,155,158,161,163,163,161,160,158,149,135,122,118,125,131,
158,158,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,159,160,160,160,160,160,159,159,159,159,160,160,160,160,159,159,160,160,160,159,159,160,159,159,159,159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,162,163,163,163,163,163,163,163,163,163,163,162,162,162,162,162,162,162,162,162,162,162,162,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,164,162,161,162,164,164,164,164,165,165,165,165,165,165,165,165,165,166,165,161,159,161,164,164,162,160,160,163,165,165,165,164,162,159,158,161,163,162,159,157,156,155,153,144,130,116,111,120,126,
159,159,159,159,159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,164,164,164,164,164,164,164,163,163,163,164,164,163,163,164,164,164,164,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,164,164,165,165,165,165,165,164,164,164,164,165,165,164,164,164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,166,166,165,165,165,165,165,165,165,165,165,166,166,165,165,166,165,161,158,160,163,164,163,163,162,163,164,165,166,166,165,166,167,167,165,158,154,157,161,161,158,157,160,164,165,166,166,166,164,161,160,163,165,165,159,153,153,155,152,142,129,118,115,120,124,
159,159,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,165,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,166,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,163,161,161,162,162,161,158,155,157,161,165,166,166,166,167,168,169,166,159,154,155,158,158,157,160,163,166,166,165,166,167,164,159,158,161,166,168,162,154,152,155,153,142,130,124,123,124,126,
160,160,160,160,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,161,162,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,165,165,165,165,165,165,166,166,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,166,166,166,166,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,167,166,163,159,157,152,148,151,158,163,164,163,163,165,168,169,167,162,156,154,156,159,161,164,167,167,166,163,162,163,161,157,155,159,165,169,164,153,149,152,152,142,131,126,127,131,133,
161,161,161,161,161,161,161,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,162,162,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,165,165,165,166,166,166,166,166,166,165,165,165,166,166,166,166,166,166,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,166,166,167,167,168,167,161,155,153,151,148,150,156,161,159,156,157,160,164,166,165,161,156,153,156,160,161,163,167,168,165,159,156,157,158,157,156,158,162,165,161,150,145,149,152,144,133,128,131,136,137,
162,162,162,162,162,162,162,162,162,162,162,163,163,163,163,162,163,163,163,162,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,162,162,162,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,163,163,163,163,164,164,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,165,166,166,166,166,166,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,167,167,167,167,166,165,164,165,165,163,159,155,154,156,157,154,153,157,159,154,149,148,150,153,157,158,157,156,155,156,156,155,157,162,165,164,160,156,156,157,159,160,160,161,162,158,148,144,149,153,148,138,135,139,139,137,
163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,163,164,164,164,164,164,163,163,164,164,164,164,164,163,164,164,164,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,168,168,167,167,166,164,163,164,164,158,149,148,155,162,164,159,156,157,158,152,143,138,136,137,143,148,152,155,154,151,149,148,149,151,155,161,164,162,160,160,162,163,163,163,162,154,144,141,145,149,146,138,138,144,143,139,
163,163,163,163,163,163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,167,167,167,167,167,167,167,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,170,170,170,169,169,169,168,166,164,164,165,167,166,160,151,150,158,165,167,162,158,159,158,150,137,129,126,129,134,138,143,150,151,148,147,145,141,138,142,155,164,163,160,160,163,164,162,162,158,147,136,133,135,138,139,136,136,140,142,142,
163,163,163,163,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,164,165,165,165,164,164,164,164,164,164,164,165,165,165,165,165,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,168,168,168,168,168,168,168,169,169,169,169,169,169,169,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,169,167,164,165,167,167,166,165,161,160,161,164,166,164,161,161,159,149,136,127,128,134,136,133,133,141,147,150,150,146,139,134,136,147,155,153,151,155,162,164,160,154,150,139,125,120,120,123,130,134,132,134,138,140,
164,164,164,164,164,164,165,165,164,164,164,165,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,166,166,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,169,166,166,166,162,160,162,164,162,159,159,161,162,160,160,158,149,137,128,132,142,142,132,126,132,142,149,151,149,147,144,140,142,144,142,144,153,162,164,156,147,142,133,120,113,112,115,123,129,129,131,136,138,
164,164,164,164,164,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,165,166,166,165,165,165,165,165,165,165,165,165,165,165,166,166,166,165,165,165,165,166,166,166,166,166,166,166,166,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,172,172,172,172,172,171,169,166,165,163,157,153,156,158,156,152,150,151,153,155,158,155,147,136,126,132,146,148,136,128,132,140,147,150,152,153,151,145,141,139,137,142,152,159,158,150,142,140,135,124,118,117,118,122,125,129,135,140,141,
165,165,165,165,165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,170,170,170,170,171,171,171,171,171,171,171,171,171,171,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,172,172,172,173,173,173,172,172,169,166,166,165,159,153,150,150,149,147,147,145,145,150,154,151,145,134,126,136,151,153,144,137,141,149,153,153,153,150,146,142,142,135,129,135,149,155,153,147,143,143,140,134,131,127,126,127,128,131,141,147,148,
165,165,165,165,165,165,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,166,167,167,167,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,173,173,173,172,172,171,171,171,172,171,165,155,148,145,147,148,149,148,146,148,148,145,143,138,134,142,152,154,148,144,152,163,164,159,151,143,138,140,144,133,119,127,147,157,156,154,150,145,141,140,137,131,128,131,132,134,142,150,152,
166,166,166,165,165,166,166,166,166,166,166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,171,171,172,172,172,172,172,172,172,172,172,172,172,173,173,173,172,171,169,170,174,178,177,169,159,151,147,147,148,152,154,150,145,141,140,143,145,143,143,147,151,152,153,162,170,166,156,145,135,133,142,147,135,120,127,147,160,164,163,157,147,141,141,138,130,126,132,136,137,141,147,149,
166,166,166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,167,168,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,168,168,169,169,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,172,172,172,173,173,173,173,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,172,173,173,172,172,171,170,165,165,171,177,175,169,162,157,152,147,146,153,158,151,142,139,140,145,148,144,139,143,152,159,165,170,169,159,148,138,132,136,146,151,144,131,131,145,161,169,168,160,152,147,146,143,135,132,138,144,144,142,141,140,
166,166,166,166,167,167,167,167,167,167,167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,169,169,169,169,169,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,172,170,170,169,164,162,167,171,172,169,166,163,157,148,146,156,162,156,147,143,145,149,148,139,132,135,147,161,171,172,166,155,144,139,141,145,150,153,149,138,133,145,163,168,164,159,155,153,151,150,148,144,146,150,149,143,139,138,
167,167,167,167,167,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,173,174,174,174,174,174,174,174,172,170,170,170,165,162,164,167,169,171,170,167,159,150,150,161,168,165,158,152,149,150,147,134,123,124,136,153,164,165,162,154,145,143,149,152,151,151,149,141,140,154,167,165,159,156,154,151,150,154,158,155,150,149,148,143,139,140,
168,168,168,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,174,174,174,175,175,175,175,175,175,173,170,170,169,165,161,161,162,164,166,165,162,156,151,154,163,168,165,160,155,149,145,140,128,119,121,134,148,155,158,158,152,142,143,152,155,152,150,150,148,152,164,170,164,159,155,149,143,144,152,161,161,153,150,151,147,140,138,
168,168,168,168,169,169,169,169,169,169,169,169,169,169,169,170,170,170,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,173,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,174,174,174,175,175,175,175,175,175,175,175,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,175,175,176,176,176,177,176,173,170,169,167,161,157,157,157,156,155,153,150,148,150,158,163,161,154,150,149,144,138,134,125,119,128,142,150,152,156,159,152,144,146,156,160,157,152,149,151,155,162,167,165,161,156,146,139,141,149,157,160,155,155,160,155,142,136,
169,169,169,169,169,169,169,169,169,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,174,174,174,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,174,170,169,167,161,154,153,153,151,148,146,143,142,149,157,159,153,145,142,144,141,137,136,128,123,135,148,150,152,160,165,163,157,157,160,161,157,147,139,141,146,154,162,164,159,154,147,143,144,147,150,153,154,158,164,159,146,140,
169,169,169,169,170,170,169,170,170,170,170,170,170,170,170,170,170,170,171,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,176,175,174,171,162,153,148,148,150,149,147,144,143,147,151,150,148,143,142,143,141,139,140,133,130,142,149,146,150,163,176,179,174,167,159,151,147,141,132,134,143,151,159,160,155,151,149,147,145,143,144,149,155,160,159,154,147,145,
170,170,170,170,170,170,170,170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,179,178,177,172,163,154,148,148,150,150,150,148,145,143,144,143,145,146,145,142,138,139,144,142,143,148,147,143,146,159,177,185,182,170,151,136,137,141,140,145,154,155,154,153,150,150,151,147,143,142,144,148,156,159,152,144,142,143,
170,170,170,170,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,171,172,172,172,172,172,172,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,176,176,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,177,172,165,160,156,153,151,150,149,152,151,143,138,141,144,148,150,147,139,135,141,152,157,157,154,147,142,144,153,167,176,175,164,142,124,130,143,150,157,164,159,148,142,144,150,151,144,138,141,147,152,158,157,148,140,142,145,
171,171,171,171,171,171,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,176,176,176,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,178,178,176,172,163,155,154,157,157,154,149,149,154,153,143,138,143,151,155,154,145,135,131,139,154,163,161,154,146,143,146,151,156,160,160,153,134,120,128,143,147,153,161,158,142,130,134,145,148,141,135,139,151,161,164,158,147,142,146,150,
171,172,172,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,174,174,173,173,174,174,174,174,174,174,174,174,174,175,175,175,174,174,175,175,175,175,175,174,174,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,178,178,178,178,179,179,179,179,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,179,179,179,175,166,156,149,152,160,161,156,152,153,158,157,148,141,146,156,159,152,138,127,122,130,144,152,152,149,143,141,146,150,149,147,149,146,134,129,137,144,141,142,149,149,134,121,125,138,144,140,136,139,152,166,169,159,147,142,144,147,
172,172,172,172,172,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,173,174,174,173,173,174,174,174,174,174,174,173,173,173,174,174,174,174,174,174,174,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,176,166,156,151,156,164,164,158,156,160,162,160,151,142,143,152,154,143,128,119,118,125,134,138,140,141,138,136,142,149,147,143,144,144,140,142,148,149,143,141,143,138,126,119,124,135,141,140,139,141,150,162,166,157,145,140,142,144,
173,173,173,173,173,173,173,173,174,174,174,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,180,175,168,162,158,161,168,164,154,154,160,162,158,151,140,136,141,145,137,125,120,124,131,133,132,134,136,134,133,141,148,147,144,142,139,139,143,148,150,148,145,142,134,124,123,127,132,135,138,141,146,152,159,159,150,141,140,145,148,
173,173,173,173,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,180,180,177,173,170,168,164,164,169,163,150,147,154,157,156,152,142,134,138,144,140,128,122,131,140,137,132,134,137,138,138,143,145,142,138,133,126,127,133,140,148,150,147,143,136,129,127,127,127,129,136,145,151,155,157,151,141,137,141,147,150,
174,174,174,174,174,174,174,174,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,181,181,181,180,180,177,175,174,172,169,170,172,170,168,170,165,152,146,151,156,157,152,144,140,145,150,145,131,122,131,141,139,136,138,144,148,148,145,138,130,128,123,117,122,131,138,146,148,145,143,139,133,128,126,125,127,136,146,149,148,146,142,138,141,144,145,145,
175,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,176,176,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,181,180,178,174,169,166,163,161,164,170,173,174,175,171,161,156,159,161,157,150,144,147,155,155,145,131,124,129,139,142,139,140,148,153,151,143,128,119,120,122,123,134,143,141,138,140,142,143,141,133,127,126,127,130,137,142,139,135,134,136,144,151,148,140,137,
175,175,175,175,175,175,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,182,181,180,180,181,179,173,165,159,154,152,155,162,169,175,176,173,168,166,165,162,155,148,144,150,156,148,136,128,125,130,140,145,141,135,136,142,141,131,117,110,115,123,132,147,155,143,129,130,138,144,141,131,123,125,131,136,142,143,136,130,132,139,151,156,146,133,130,
176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,176,176,177,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,181,174,170,174,181,181,175,163,152,149,151,155,158,161,165,166,165,163,162,161,158,154,150,146,145,141,131,122,121,124,131,140,146,141,127,120,124,124,116,108,109,117,123,129,145,156,143,126,125,134,138,136,126,119,124,137,148,155,152,141,133,134,139,147,150,138,125,122,
176,176,176,176,176,176,176,176,176,176,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,183,182,183,182,181,178,168,161,168,179,182,175,161,149,151,160,163,158,151,152,154,155,154,154,155,157,158,157,153,142,130,119,115,117,123,130,137,144,143,128,115,114,114,112,112,121,132,130,123,130,143,141,131,129,130,129,127,122,117,125,142,159,166,159,145,134,129,129,133,136,130,119,114,
177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,187,186,181,178,181,182,180,177,170,165,170,177,177,170,157,150,159,169,167,154,145,148,155,157,157,156,157,161,163,164,161,149,134,124,121,121,122,126,133,143,146,133,115,112,117,120,123,134,144,138,122,120,130,136,139,139,133,128,125,120,116,124,143,160,166,157,142,131,126,123,123,128,127,118,113,
177,177,177,177,177,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,183,183,184,184,184,184,184,184,184,184,184,184,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,187,189,185,174,170,176,180,179,178,178,176,177,176,171,162,152,152,163,169,161,147,144,154,163,166,163,160,159,162,163,162,159,152,142,135,132,128,123,123,131,142,145,130,111,112,124,128,130,137,142,135,123,118,121,128,136,141,139,136,132,125,120,127,144,156,156,146,133,127,128,128,125,127,130,127,123,
178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,178,179,178,178,179,179,179,179,178,178,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,183,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,184,185,185,185,185,185,184,184,185,185,185,185,185,185,184,185,185,185,185,185,185,185,185,187,190,189,177,162,162,171,176,174,174,177,179,179,176,170,161,152,152,160,160,149,142,146,160,170,168,160,154,155,159,159,154,149,144,139,138,138,133,126,126,131,138,135,120,108,116,131,131,126,129,132,127,121,120,122,125,130,134,139,143,141,134,130,136,148,152,144,133,124,121,125,128,124,124,130,133,133,
179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,188,191,183,162,151,159,170,170,165,163,167,172,174,172,170,163,155,153,152,149,142,141,150,164,169,161,148,142,147,154,154,147,141,135,130,131,135,132,126,126,129,132,126,112,110,125,137,131,122,121,124,121,119,125,132,134,131,129,135,145,143,135,132,139,148,148,141,132,125,121,119,118,116,116,121,130,134,
179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,185,168,148,147,163,171,164,155,153,158,163,165,166,167,163,155,147,141,138,139,145,155,163,161,151,139,135,140,147,148,143,136,131,126,123,124,123,121,121,124,127,121,111,116,133,140,131,120,118,121,124,127,136,146,144,136,130,135,141,134,121,121,133,142,145,146,144,140,134,123,116,116,114,116,130,138,
179,179,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,186,178,157,141,150,169,173,162,153,153,158,162,162,163,164,160,149,137,130,131,139,150,157,156,151,144,139,136,138,142,144,141,134,132,132,125,116,113,115,118,120,120,115,112,122,137,138,127,119,118,126,135,142,149,152,146,138,135,136,134,119,105,110,127,138,144,150,152,151,147,137,132,129,120,119,135,146,
180,180,180,180,180,181,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,180,180,180,180,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,187,178,160,146,155,172,174,165,157,158,163,164,164,164,162,156,146,135,131,134,143,152,154,150,145,140,139,138,137,138,141,142,138,139,141,132,117,114,121,126,125,117,111,115,130,142,138,127,122,124,134,145,149,150,150,144,142,143,141,132,112,97,103,121,134,143,150,150,145,145,149,150,140,122,119,137,149,
181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,183,168,154,159,173,177,172,165,162,165,165,164,165,163,159,154,148,144,144,146,148,152,153,148,139,136,139,139,135,137,143,143,142,140,131,123,127,138,140,132,120,113,119,137,149,146,136,131,132,139,145,143,140,142,145,149,151,147,138,119,99,99,116,133,145,151,145,135,138,153,157,140,119,117,135,146,
181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,182,181,181,181,181,181,181,181,181,181,181,181,181,182,182,182,182,182,182,182,182,182,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,186,186,186,187,187,187,187,187,187,187,186,186,186,187,187,187,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,188,183,168,156,161,174,179,176,171,167,166,164,163,165,166,166,164,160,155,151,147,145,152,159,155,145,141,145,145,137,131,134,138,137,131,124,127,141,152,146,131,118,114,123,140,153,150,140,136,138,139,138,133,131,137,147,152,153,153,150,135,113,107,122,140,150,151,140,129,133,149,154,141,126,123,134,142,
182,182,182,182,183,183,182,183,183,183,183,183,183,183,183,183,183,183,183,182,182,182,182,182,182,182,182,182,182,181,182,182,182,182,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,188,181,167,157,163,174,178,176,172,168,164,162,162,163,165,166,166,162,158,154,149,146,151,157,156,150,148,149,147,138,125,121,126,131,129,126,133,149,156,144,127,116,116,127,139,144,138,130,132,140,140,130,123,125,136,146,148,149,155,155,141,123,119,130,143,151,149,138,129,132,143,150,149,139,132,135,139,
182,182,183,183,183,183,183,183,183,183,183,184,183,183,183,184,184,183,183,183,183,183,183,182,182,182,182,182,182,182,182,182,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,187,188,188,188,188,188,188,188,188,188,188,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,182,170,163,167,173,173,171,168,162,160,162,163,164,165,165,162,159,158,156,151,148,150,151,150,148,146,142,140,135,125,117,119,127,133,136,142,153,157,147,130,120,121,128,131,125,119,119,128,140,142,127,113,117,130,138,136,138,145,143,130,122,121,126,133,141,144,141,138,137,140,149,152,142,133,133,136,
182,183,183,183,183,183,183,183,183,184,184,184,184,184,184,184,184,184,184,184,183,183,183,183,183,182,182,182,182,182,183,183,183,184,184,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,187,187,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,191,190,185,178,171,171,172,171,168,163,156,157,163,167,168,169,168,163,158,157,156,151,149,148,147,146,145,141,137,135,134,129,121,119,127,137,145,150,153,155,151,136,120,120,126,126,117,111,116,127,139,141,127,110,110,118,122,120,122,130,130,125,122,122,120,125,135,142,147,151,146,137,138,141,134,127,129,131,
175,176,176,177,177,177,177,178,177,177,177,178,178,178,177,179,179,179,179,179,178,179,179,178,179,180,180,179,180,182,183,183,184,184,184,185,185,185,185,185,185,185,185,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,191,190,187,180,174,172,171,169,163,158,160,166,171,174,174,171,165,159,155,151,148,147,147,147,145,141,137,139,139,135,128,121,120,129,141,152,155,150,146,145,133,118,118,129,134,128,123,124,129,135,137,130,122,117,110,105,105,114,124,130,131,129,124,122,130,141,146,153,158,146,123,116,122,127,126,125,125,
146,147,148,151,152,152,154,155,154,153,153,155,156,154,155,160,161,160,162,161,159,162,161,157,160,165,164,164,172,180,183,184,184,184,185,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,187,187,188,188,188,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,189,189,189,190,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,192,192,192,192,191,191,192,192,192,192,192,192,192,192,192,192,192,192,194,198,196,185,175,173,173,170,165,162,164,168,174,176,175,171,166,159,150,145,146,147,147,148,143,133,131,139,139,128,118,114,115,125,139,151,153,143,132,130,126,121,126,136,142,141,140,140,136,132,132,134,135,128,112,101,103,112,121,128,131,128,123,128,141,149,149,152,152,134,107,100,113,127,128,124,122,
98,98,100,104,109,114,119,123,123,121,122,123,124,123,126,132,133,132,134,132,130,134,131,122,124,129,127,133,156,177,183,183,184,185,185,185,186,186,186,186,186,186,186,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,188,188,188,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,193,193,193,193,194,199,205,198,177,162,162,166,166,163,162,164,170,175,174,170,166,164,157,147,144,148,150,150,150,143,131,130,137,134,120,113,111,109,112,124,139,145,136,124,118,116,122,132,138,138,141,149,153,148,136,131,135,138,131,120,115,115,114,115,120,125,125,126,134,144,145,142,145,142,122,101,99,114,127,128,121,117,
61,61,62,68,76,86,96,104,105,105,106,106,106,105,107,111,112,112,114,111,108,111,106,94,89,87,86,104,142,173,183,183,184,185,185,186,186,186,186,186,186,187,187,187,187,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,189,189,189,189,188,189,189,189,189,189,189,189,189,190,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,190,190,190,190,190,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,194,197,205,209,191,158,136,136,146,155,159,163,168,172,174,169,161,159,162,158,150,148,152,154,154,154,148,138,136,136,129,121,120,118,108,104,113,130,139,135,125,114,108,115,129,135,133,137,150,159,155,144,138,140,139,132,131,133,129,119,112,113,119,127,131,136,137,133,132,139,138,121,105,106,114,119,119,114,110,
58,58,59,64,72,81,91,98,101,104,103,102,102,101,101,104,104,103,106,106,101,98,94,84,73,63,62,85,131,168,182,184,184,185,186,186,186,187,187,187,187,187,187,187,187,187,187,188,188,188,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,191,191,191,191,191,191,191,191,191,191,190,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,191,191,191,191,191,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,194,194,194,194,194,194,194,194,194,194,194,194,194,195,200,209,211,190,152,123,117,128,146,159,169,177,178,176,167,155,153,159,162,158,154,155,156,157,155,149,144,142,135,128,129,136,132,117,107,113,127,135,134,127,115,106,113,129,136,134,138,151,158,157,155,153,149,144,139,139,140,133,122,113,110,112,120,125,127,126,123,127,137,137,122,111,112,112,109,112,115,114,
75,75,76,78,80,84,92,97,100,102,99,98,100,98,95,98,98,96,100,105,100,94,88,78,65,53,49,67,113,157,179,184,185,185,186,186,187,187,187,188,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,192,192,191,191,191,191,191,191,191,191,191,191,190,190,190,190,189,189,189,189,189,189,189,189,189,189,189,189,189,190,190,191,191,191,191,192,192,192,192,192,193,193,193,193,193,193,194,194,194,194,194,194,194,194,195,195,195,195,195,195,195,195,195,195,195,195,198,203,212,216,201,168,138,126,131,148,164,177,183,183,179,170,154,148,155,161,162,159,156,158,159,152,144,143,143,138,133,141,152,150,133,117,113,118,123,123,117,110,109,124,144,149,139,137,146,152,155,161,157,145,139,141,143,140,130,121,116,111,106,106,113,118,116,114,121,132,132,121,116,120,115,107,115,126,129,
90,89,88,88,86,86,92,97,100,100,97,95,97,95,90,92,94,91,94,103,102,92,81,69,56,43,35,47,91,145,176,184,185,186,186,187,187,188,188,188,188,188,188,188,188,189,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,192,192,192,192,192,192,192,192,192,191,191,191,191,191,190,190,189,189,189,189,189,189,188,188,188,189,189,189,189,190,190,191,191,191,192,192,192,192,193,193,193,194,194,194,194,194,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,196,197,200,206,217,225,214,185,161,150,151,160,171,178,181,182,180,171,155,148,153,159,164,164,159,158,158,150,142,143,147,145,142,148,157,160,150,129,112,105,105,105,103,105,119,142,162,159,138,129,133,138,144,149,139,123,121,132,141,139,129,121,119,115,106,102,111,119,115,109,116,128,130,125,126,130,123,116,124,136,139,
97,95,91,89,89,88,92,99,101,99,99,98,97,95,91,91,93,91,92,99,98,84,68,56,45,31,23,34,78,136,173,184,185,186,187,187,188,188,189,189,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,192,189,187,186,185,185,187,189,191,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,193,192,192,192,192,192,192,191,191,191,190,190,189,189,189,188,188,188,188,188,188,189,189,189,190,190,191,191,192,192,192,192,193,193,194,194,194,194,194,195,195,195,195,195,195,195,195,195,195,195,195,195,195,196,196,196,196,196,196,197,201,206,213,226,234,221,192,172,166,166,170,172,172,173,175,175,168,156,150,154,160,166,166,160,154,151,146,144,148,154,153,148,147,152,158,159,143,117,99,93,93,98,111,133,158,169,154,131,125,128,127,127,127,116,101,102,117,133,138,133,125,122,117,109,107,116,125,121,115,122,133,133,127,128,132,129,129,136,142,143,
96,93,88,89,91,89,92,98,98,97,101,101,97,94,92,91,91,88,90,93,88,71,57,47,35,22,17,29,69,125,167,182,185,186,187,188,188,189,189,189,190,190,190,190,190,190,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,193,193,191,184,174,167,163,163,170,182,190,192,193,193,193,193,193,193,193,194,194,194,194,194,194,194,194,194,194,194,194,194,194,193,193,193,193,193,193,193,192,192,192,191,191,190,190,189,189,188,188,187,185,184,185,187,188,189,189,190,190,191,191,192,193,193,193,193,194,194,195,195,195,195,195,195,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,196,197,201,209,216,222,233,239,223,194,175,170,171,172,166,160,163,168,168,162,155,151,153,158,164,165,159,150,144,143,147,152,157,156,149,145,144,150,158,148,124,106,99,99,102,112,134,159,165,147,130,128,128,121,115,115,109,96,92,104,120,131,134,132,126,118,112,112,119,126,125,123,129,137,130,115,111,117,124,132,142,147,147,
93,90,88,92,92,89,91,96,95,95,101,101,94,89,91,93,90,86,86,88,80,65,53,42,27,17,14,24,55,106,154,179,185,187,188,188,189,189,190,190,190,191,191,191,191,191,191,191,191,191,191,191,192,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,192,193,193,193,193,193,194,194,193,193,193,193,193,194,194,191,179,161,145,135,133,145,170,188,193,193,193,193,194,194,194,194,194,194,194,194,195,194,194,194,194,194,194,194,194,194,194,194,194,194,194,194,193,193,193,192,192,191,191,190,189,188,188,187,181,170,163,171,182,188,189,189,190,190,191,192,192,193,193,194,194,194,195,195,195,195,195,196,196,196,196,196,196,196,196,197,197,197,197,196,196,196,197,197,197,197,198,206,219,225,224,230,236,222,194,175,170,171,169,158,149,153,161,162,159,156,153,151,153,160,164,161,152,147,149,154,156,157,154,148,140,134,137,145,141,126,120,118,115,109,105,118,146,158,145,129,126,123,114,110,114,113,103,95,102,114,122,129,135,130,120,114,117,123,127,128,127,131,132,118,100,92,96,105,116,130,141,145,
97,93,92,95,95,90,92,96,97,98,100,101,95,89,93,99,98,92,86,81,74,68,58,40,22,14,13,18,40,88,144,177,186,187,188,189,190,190,190,191,191,191,191,191,191,192,192,192,192,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,193,193,193,194,194,194,194,194,194,194,194,194,194,194,194,194,192,181,162,143,130,124,135,164,186,193,193,193,194,194,194,194,194,194,194,195,195,195,195,195,195,195,195,195,195,195,195,194,194,194,194,194,194,194,193,193,193,192,192,191,190,189,188,187,181,163,134,120,137,167,183,188,189,190,191,191,192,193,193,194,194,194,195,195,196,196,196,196,196,196,197,197,197,197,197,197,197,197,197,197,197,197,197,197,198,198,198,201,212,226,227,216,216,227,220,193,174,170,171,167,155,144,144,154,160,159,158,157,153,153,159,163,161,157,156,158,159,158,155,154,149,138,128,129,135,132,126,126,127,123,113,100,103,127,150,145,127,120,118,112,112,117,114,107,106,115,121,120,125,132,128,116,113,123,132,132,130,132,133,127,111,94,88,90,93,98,111,128,136,
107,102,96,97,98,95,93,97,101,102,100,102,100,94,94,102,108,102,85,69,65,71,69,46,22,14,13,16,34,80,138,174,185,187,189,190,190,190,191,191,191,191,192,192,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,193,194,194,194,194,194,194,194,193,194,194,194,194,194,194,194,194,194,194,194,194,194,193,186,174,161,149,138,141,164,186,193,193,193,194,194,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,195,194,194,194,194,193,193,192,191,190,189,188,182,163,127,86,71,94,135,168,184,189,190,191,192,192,193,194,194,195,195,195,196,196,196,196,197,197,197,197,197,197,197,198,198,198,198,198,198,198,198,198,198,200,200,200,204,216,225,217,199,199,216,217,193,174,170,173,171,162,151,147,152,160,161,159,160,162,163,164,163,162,163,163,162,158,155,156,159,153,141,134,133,132,127,121,121,123,125,122,111,100,112,137,142,125,114,113,113,117,116,109,107,115,128,132,127,128,132,124,110,111,127,140,136,131,135,135,126,110,97,96,102,101,98,109,125,131,
111,105,97,96,98,96,94,98,103,103,101,103,103,97,94,102,110,103,80,61,61,77,83,61,30,15,12,14,29,67,122,165,183,188,189,190,191,191,191,191,192,192,192,192,192,192,193,192,193,193,193,193,193,193,193,193,193,193,193,193,193,193,194,194,194,194,194,194,194,193,194,194,194,194,194,195,195,194,193,191,191,191,191,191,188,181,175,166,149,142,157,176,183,184,186,189,192,193,194,195,195,195,195,196,196,196,196,196,196,196,196,196,196,196,196,196,195,195,195,195,194,194,194,194,193,192,192,191,189,183,164,128,83,49,40,58,94,136,168,185,190,192,192,193,194,194,195,195,195,196,196,197,197,197,197,197,198,198,198,198,198,198,198,199,199,199,199,199,199,199,200,201,202,201,206,218,218,201,182,186,210,215,192,174,171,176,177,173,165,161,161,162,161,160,164,169,170,165,160,162,167,168,164,157,152,155,162,158,151,148,143,132,121,116,118,124,131,138,131,109,100,114,124,117,107,104,109,117,114,109,112,122,130,135,138,140,139,129,116,116,128,136,131,129,136,139,129,112,98,100,113,115,111,121,134,139,
104,102,99,97,97,97,97,100,103,103,103,104,102,96,96,103,103,88,68,58,66,86,99,79,41,17,12,13,21,48,97,150,180,188,189,190,191,191,192,192,192,192,192,192,193,193,193,193,193,193,193,193,193,194,194,194,194,194,194,193,193,193,194,195,195,195,195,195,194,194,194,195,195,195,195,195,195,192,185,179,177,176,175,180,184,182,177,168,144,122,124,137,145,150,157,168,179,184,185,187,190,191,191,191,190,190,190,192,192,193,193,194,193,193,192,192,192,192,192,191,190,189,189,188,188,188,188,188,182,164,128,83,47,30,28,38,59,94,136,169,184,188,190,191,192,193,195,195,196,196,197,197,197,197,198,198,199,199,199,199,199,199,199,199,200,200,200,200,199,199,200,201,201,199,206,217,210,188,173,183,209,215,192,174,172,177,179,176,174,173,168,163,159,160,165,168,165,157,151,154,164,168,164,157,150,150,156,160,163,163,152,135,123,120,123,127,132,142,142,122,100,94,98,103,103,101,110,123,121,119,126,128,124,131,145,152,149,142,134,129,128,125,120,124,137,143,131,110,96,99,111,117,117,128,141,146,
95,98,100,99,98,98,100,101,100,101,104,105,100,96,98,102,93,73,59,60,74,95,109,93,52,21,12,12,15,34,80,139,177,188,189,190,191,191,192,192,192,193,193,193,193,193,193,193,194,194,194,194,194,194,194,195,195,195,194,194,194,194,195,195,196,195,195,195,195,195,195,195,196,196,196,196,194,187,171,158,156,154,151,159,170,171,167,156,126,91,78,85,91,97,108,126,147,161,164,166,171,176,177,173,168,166,168,171,174,177,179,181,181,181,178,176,176,175,175,174,171,168,165,164,166,169,172,171,157,124,81,46,28,22,22,26,38,60,96,135,162,173,179,182,184,187,189,190,191,192,193,193,192,193,193,193,194,194,194,195,195,195,196,196,197,196,196,196,196,195,196,197,195,194,199,205,198,180,170,185,212,216,193,175,173,176,174,171,172,172,166,161,159,161,163,159,151,143,138,141,152,159,157,151,145,142,145,155,167,169,157,142,134,130,126,123,121,129,137,130,111,95,90,95,103,108,119,132,133,136,143,136,121,123,140,152,154,153,150,141,130,120,114,118,133,140,126,108,103,107,112,114,115,126,140,144,
90,94,98,99,98,98,100,98,94,96,101,104,100,96,97,95,83,66,61,70,84,99,111,101,64,28,13,11,13,27,68,126,169,186,190,191,191,192,192,193,193,193,193,194,194,194,194,194,194,194,195,195,195,195,195,195,195,195,194,194,195,195,196,196,196,196,196,196,196,196,196,196,197,197,197,196,191,175,149,134,135,137,135,136,140,140,138,131,106,71,59,66,68,68,76,90,110,128,133,133,139,149,151,143,134,131,135,142,147,152,155,157,161,160,154,152,151,150,150,146,139,134,130,130,133,138,141,136,113,76,44,27,21,19,17,19,28,41,63,94,126,149,162,168,170,172,171,170,171,172,174,174,173,174,173,173,175,175,173,177,179,180,181,182,183,182,181,181,181,180,181,180,176,175,177,179,175,166,165,188,218,219,194,177,174,172,165,160,162,163,159,160,163,162,158,150,139,131,129,134,143,147,145,142,140,138,139,147,157,161,153,145,140,132,122,115,114,121,130,131,124,116,108,102,103,113,127,137,140,148,155,147,128,120,130,142,146,150,155,148,132,120,112,114,122,127,119,113,120,126,124,117,115,124,134,136,
87,89,93,94,94,97,98,95,90,90,96,99,97,94,91,84,71,63,69,82,92,99,109,108,79,39,16,10,12,21,52,105,156,183,190,191,192,192,193,193,193,194,194,194,195,195,195,195,195,195,195,196,196,196,196,196,196,195,194,193,194,195,196,197,197,196,196,197,197,196,196,196,197,198,197,196,188,161,125,111,121,130,128,118,110,108,109,109,96,75,74,86,85,78,80,86,96,106,110,110,116,127,131,124,113,113,120,125,132,139,138,139,145,144,138,138,139,139,140,134,124,118,114,113,118,118,110,93,67,40,26,21,19,18,16,17,22,32,45,63,91,122,145,154,155,153,146,138,134,134,140,145,146,148,149,149,153,153,150,154,160,161,162,163,164,162,160,160,160,158,157,153,149,151,152,153,153,152,164,196,225,220,194,177,174,169,156,146,148,152,153,160,165,159,148,142,138,135,135,139,141,140,139,142,146,144,140,141,146,148,144,138,134,127,115,108,114,125,131,131,131,136,135,117,105,117,134,139,141,151,162,159,144,131,131,134,133,141,154,150,133,117,108,107,109,111,113,120,132,138,133,124,118,122,127,126,
83,84,87,90,92,94,96,95,90,87,89,89,88,88,83,71,61,63,77,90,96,99,107,112,90,48,19,12,12,17,38,87,145,181,190,192,192,193,193,194,194,194,195,195,195,196,196,196,196,196,196,196,196,196,197,197,197,196,194,192,192,194,196,197,197,196,196,197,197,196,196,196,197,197,197,195,185,155,117,102,113,123,121,110,100,98,101,103,100,93,96,110,111,103,102,106,109,109,110,114,119,126,132,127,115,117,125,127,133,141,136,134,142,140,135,141,144,145,150,144,134,131,126,122,124,115,87,57,36,24,19,19,19,19,18,18,20,25,35,47,65,92,121,137,139,136,129,116,106,107,117,129,134,140,145,147,152,154,150,152,157,158,159,159,157,155,153,154,153,150,145,142,141,145,148,150,153,159,178,211,233,221,192,176,174,169,151,134,135,143,150,159,162,150,137,136,144,149,148,145,142,141,142,148,155,154,144,140,143,143,137,129,126,123,113,104,112,129,135,130,128,142,150,133,114,120,134,137,138,151,166,169,159,147,141,136,127,134,149,149,131,112,102,103,103,103,109,121,130,130,128,123,118,118,116,114,
84,85,88,91,91,91,93,96,93,87,83,79,79,81,75,63,60,71,85,95,98,98,104,109,93,55,25,16,15,17,33,77,135,176,189,192,193,193,194,194,195,195,195,196,196,196,196,196,196,197,197,197,197,197,197,197,197,197,195,192,191,193,196,197,197,196,196,197,197,197,197,197,197,196,195,193,180,151,121,107,112,119,118,112,108,107,105,107,112,113,118,129,132,124,122,128,127,121,124,130,133,139,146,138,124,125,131,131,138,144,136,133,141,137,133,144,148,149,156,154,146,146,138,124,118,100,64,34,22,18,17,18,19,20,20,20,19,21,27,37,48,65,89,110,118,123,128,122,114,116,126,138,145,152,159,162,165,168,166,165,167,167,166,166,163,161,162,163,162,160,156,154,157,160,163,167,172,181,200,226,238,220,190,175,175,171,151,129,128,140,151,160,160,146,135,136,147,154,152,148,146,144,145,150,159,161,151,144,147,145,134,126,125,125,114,101,106,125,134,125,121,136,150,138,119,116,124,129,135,151,169,176,169,154,145,137,126,126,137,139,125,107,101,108,111,105,102,108,114,110,106,106,106,105,102,98,
97,96,94,95,95,94,96,96,93,89,87,85,84,83,72,62,67,81,93,98,99,98,101,105,92,59,30,20,18,19,31,65,119,165,187,192,193,194,194,195,195,196,196,196,196,197,197,197,197,197,197,197,197,198,198,198,197,196,195,194,194,195,196,198,198,197,196,196,197,198,198,197,196,195,194,189,168,137,116,112,118,124,122,119,120,117,112,118,128,133,139,146,143,134,134,137,129,124,129,133,133,142,149,138,127,129,130,128,135,139,131,130,134,128,127,136,139,139,145,144,140,142,131,106,84,63,39,24,18,16,16,18,20,21,22,21,20,18,21,28,38,49,63,80,96,115,134,142,142,145,150,152,154,159,162,163,166,170,169,167,167,165,164,163,162,163,164,165,166,168,166,165,168,170,172,178,184,193,210,232,240,220,190,176,175,167,143,120,121,140,155,164,164,154,146,145,150,153,152,152,150,141,135,141,153,162,159,154,152,143,131,128,133,129,115,104,108,122,127,117,113,126,138,132,117,107,110,120,130,148,170,181,174,159,146,137,126,120,123,126,120,108,107,119,123,106,90,91,100,99,90,86,88,88,85,84,
108,104,97,95,100,106,104,95,88,89,94,97,94,86,73,67,76,89,97,99,99,98,99,102,92,63,35,23,20,21,27,51,99,153,184,192,193,194,195,195,196,196,196,197,197,197,197,198,198,198,198,198,197,197,198,198,197,195,194,195,196,197,198,199,199,198,196,195,196,199,199,197,196,196,195,186,156,120,105,111,124,128,125,125,127,122,122,132,138,138,143,145,135,128,131,128,120,119,124,123,123,131,136,130,126,127,125,125,130,130,129,130,129,126,128,131,132,133,133,130,130,131,116,84,52,32,23,20,18,17,17,19,21,22,22,22,20,18,18,21,30,40,50,61,80,108,135,152,157,157,154,149,146,149,150,149,154,158,157,156,155,150,150,152,152,155,157,157,160,165,164,161,162,162,164,170,177,187,208,232,240,222,193,178,173,153,120,97,102,129,154,168,172,169,163,157,155,157,158,155,147,130,120,129,143,152,156,157,150,134,124,130,139,134,120,118,125,125,116,110,113,122,128,124,111,97,98,111,122,138,162,178,174,162,149,142,135,126,123,129,130,121,117,130,133,112,91,93,105,108,97,89,86,83,81,82,
109,105,96,93,101,111,108,94,85,86,91,92,86,76,70,74,85,94,98,100,100,99,99,100,93,73,47,28,20,20,23,39,83,142,180,192,194,195,195,196,196,197,197,197,197,198,198,198,198,199,199,199,198,197,197,197,197,195,194,195,197,198,200,200,200,198,194,191,195,199,200,198,197,198,196,181,149,117,105,113,125,127,124,127,128,124,127,134,130,125,127,126,118,115,118,117,116,117,117,117,120,124,129,133,133,129,130,134,131,131,138,139,134,137,141,137,138,144,141,135,137,134,112,77,43,23,17,18,18,18,19,20,21,22,22,22,21,19,18,19,24,31,39,50,68,95,125,147,153,149,143,140,139,140,143,146,150,154,154,154,152,147,146,150,153,156,159,159,163,168,167,162,158,154,154,161,168,178,203,231,240,224,196,180,169,137,91,63,69,104,144,168,177,179,174,165,159,158,154,146,135,121,118,130,140,141,142,144,137,124,119,127,136,132,125,134,144,133,111,107,121,133,133,122,104,91,97,111,119,130,150,166,166,157,151,152,150,140,135,144,144,127,118,132,139,125,113,116,123,125,119,113,107,100,97,97,
105,103,99,95,98,103,99,92,91,93,90,80,68,60,64,77,90,97,99,100,100,100,99,99,99,91,67,37,20,17,18,30,67,124,170,190,194,195,196,196,197,197,197,198,198,198,199,199,199,199,199,199,199,197,196,196,196,195,194,194,194,196,199,200,200,198,191,188,192,198,200,200,199,199,193,171,140,121,116,119,126,128,128,131,131,126,127,127,120,112,113,117,116,113,116,122,123,117,115,123,128,126,132,143,142,135,141,145,136,135,147,145,138,146,150,141,143,156,153,145,147,143,119,85,50,25,14,15,18,20,21,20,21,21,22,22,21,22,22,21,20,20,26,37,55,85,119,142,151,150,146,148,148,146,149,154,155,158,161,159,155,152,151,153,159,166,169,169,173,177,177,173,166,157,155,164,173,183,205,231,241,225,198,180,166,129,75,41,43,78,128,162,175,177,173,167,160,152,142,133,124,121,129,140,142,134,128,128,124,118,118,127,130,124,124,139,153,141,114,107,127,144,142,128,109,99,107,121,127,129,139,153,159,156,157,163,163,151,142,143,137,117,110,124,132,129,131,137,139,139,137,137,133,126,119,117,
100,101,101,99,94,89,87,91,101,107,97,78,62,55,63,80,93,98,99,100,101,100,99,99,104,105,84,47,21,14,14,21,48,100,156,187,194,195,196,196,197,198,198,198,199,199,199,200,200,200,200,200,200,198,197,197,196,194,193,192,190,190,195,199,200,198,192,187,190,195,198,200,200,198,187,158,127,118,122,124,129,133,137,140,137,131,129,127,118,113,119,128,126,122,126,131,125,113,117,130,131,125,129,138,136,132,141,144,134,133,142,138,133,144,146,135,139,152,150,141,142,139,120,94,61,29,13,13,18,22,23,22,20,20,21,22,23,26,30,28,21,14,14,24,45,83,125,148,156,160,158,156,156,153,150,150,151,153,155,153,148,147,147,147,154,166,169,166,167,172,175,174,167,160,161,171,181,192,208,228,238,225,198,179,165,129,74,37,33,58,106,151,169,166,160,159,158,150,140,131,123,125,137,144,138,129,122,120,118,115,118,125,126,120,122,139,157,151,123,108,123,141,142,133,120,111,115,127,134,133,134,145,158,166,169,171,169,156,139,129,119,109,111,122,122,119,129,142,146,143,141,142,142,139,132,128,
95,96,98,98,93,87,85,91,101,103,91,74,63,62,72,85,95,99,100,101,101,101,100,100,104,108,95,59,27,14,13,16,35,83,144,183,194,195,196,197,198,198,199,199,199,200,200,200,201,201,201,201,201,199,198,198,196,191,188,190,189,189,194,199,201,199,193,188,189,191,193,196,197,193,177,145,117,111,118,123,128,134,142,142,135,132,132,128,119,118,128,133,128,126,130,129,118,111,118,128,128,121,120,124,126,128,133,136,133,133,132,129,131,139,136,129,135,143,138,132,134,129,113,94,65,31,13,13,20,25,26,24,22,23,24,24,26,32,41,39,26,12,8,15,39,81,126,150,155,155,150,145,145,146,140,136,139,144,146,145,145,147,146,144,150,161,161,156,157,162,168,169,162,158,165,172,178,187,198,214,227,221,197,179,167,131,75,36,28,42,82,132,160,157,149,151,154,151,145,135,125,130,143,147,139,129,121,115,112,111,114,119,120,120,128,146,163,162,136,113,120,137,140,132,124,118,117,126,139,144,140,140,153,170,175,173,167,154,133,116,110,114,125,131,122,110,118,136,142,138,135,139,142,139,135,133,
95,94,92,92,92,91,89,88,86,81,72,64,64,72,83,93,98,101,101,102,102,102,101,99,101,107,104,76,38,17,13,15,28,69,129,174,192,196,197,198,198,199,199,200,200,200,201,201,201,201,201,202,201,199,198,199,197,191,187,191,192,192,195,199,201,199,194,189,188,188,189,193,193,183,162,131,110,109,116,122,126,135,143,136,125,125,130,127,119,118,124,126,123,124,128,129,123,116,115,121,127,124,119,123,133,133,127,131,141,142,132,130,140,142,131,130,142,144,133,132,139,131,108,84,57,28,13,15,22,27,28,26,27,29,29,27,28,36,48,47,30,13,6,11,33,72,114,143,151,145,136,135,138,139,136,135,140,148,151,154,160,163,160,156,160,164,161,157,159,165,171,174,168,164,171,177,179,182,186,195,211,213,195,180,167,130,73,34,26,33,61,107,143,152,149,149,150,150,148,138,127,133,149,156,150,137,121,109,105,108,114,114,114,122,138,155,166,163,140,120,127,142,141,129,124,127,130,136,148,155,150,139,140,156,169,171,165,149,124,108,112,126,138,138,123,111,116,130,134,131,134,145,148,140,133,132,
100,96,90,87,86,86,87,82,71,62,60,61,69,83,93,98,100,102,103,103,103,102,101,99,99,106,110,89,50,22,14,14,23,53,107,160,189,196,197,198,199,199,200,200,200,201,201,201,201,202,202,202,201,199,198,199,199,194,191,193,193,190,190,195,199,200,196,191,188,186,189,193,190,175,146,116,103,109,120,125,130,141,147,134,118,120,131,131,121,115,118,123,123,124,132,142,137,121,112,121,130,125,122,132,143,136,123,129,148,150,135,134,147,146,132,134,150,148,133,135,148,136,102,72,49,27,18,22,26,27,27,26,30,33,32,28,28,37,50,49,32,14,6,9,27,58,96,132,151,147,139,143,147,141,137,143,150,155,158,163,169,169,164,161,162,160,155,154,159,165,172,176,173,168,173,184,188,189,186,186,196,200,187,172,157,118,65,33,28,31,46,80,123,148,154,153,151,152,153,145,136,138,150,158,155,141,123,111,110,116,122,121,120,128,144,158,162,152,133,126,137,147,142,132,131,141,147,149,153,158,156,143,130,135,154,169,167,142,112,103,117,132,138,132,118,113,119,123,120,120,133,150,152,139,127,124,
101,98,94,92,90,87,86,79,64,53,55,66,80,92,98,101,102,104,105,105,104,103,101,99,99,103,109,98,63,30,16,14,18,38,88,149,186,196,198,198,199,200,200,201,201,201,202,202,202,202,202,202,201,200,199,199,200,198,195,194,191,185,185,191,197,200,199,193,187,186,192,194,188,170,139,109,102,113,123,127,133,146,149,132,118,124,138,136,122,116,122,127,122,121,134,145,135,117,114,126,132,126,125,134,138,128,121,132,147,143,130,132,144,142,131,135,148,142,127,133,146,131,97,76,65,47,33,32,31,27,24,24,27,29,29,26,27,36,49,48,31,14,7,8,20,42,72,107,136,146,144,146,145,137,133,142,152,152,151,155,158,154,151,154,157,151,146,147,152,155,160,167,166,161,165,178,186,189,190,186,184,182,169,152,134,99,57,37,35,37,42,66,107,141,154,158,159,163,163,156,149,147,149,151,149,139,129,126,127,131,137,139,139,141,147,154,154,142,131,133,144,148,146,144,145,147,145,141,145,155,162,155,136,126,141,165,165,136,111,108,118,125,126,121,111,109,113,111,106,107,121,139,142,130,118,114,
96,97,101,105,104,99,93,81,61,50,55,72,87,96,100,105,110,111,109,106,104,103,102,100,98,100,107,106,79,41,19,14,15,31,76,138,182,196,198,199,200,200,201,201,201,202,202,202,203,203,202,202,201,199,198,198,199,199,197,195,192,188,187,192,198,202,202,193,185,186,193,194,183,160,131,112,110,119,128,128,130,140,142,131,123,129,137,134,126,123,125,124,119,122,131,132,123,119,125,135,138,137,136,132,123,118,128,142,141,129,126,138,143,134,127,137,144,132,122,136,148,130,103,100,107,89,59,44,36,27,22,21,22,23,24,24,25,32,42,42,28,14,8,8,15,28,47,71,101,124,136,137,131,127,132,144,152,150,145,146,145,143,145,154,160,156,150,151,152,152,154,160,162,160,162,170,176,182,189,186,177,168,150,130,113,88,62,55,61,65,66,77,103,132,150,161,172,178,172,160,154,152,151,150,148,141,137,140,143,147,155,158,155,151,146,142,142,141,139,142,148,152,155,158,156,145,128,121,132,153,168,171,158,140,140,156,160,143,128,124,117,110,109,109,105,103,101,99,98,99,107,122,125,116,109,107,
92,95,100,104,104,102,96,81,61,54,64,81,93,98,102,111,121,122,115,109,106,104,103,101,99,99,106,110,90,51,22,13,13,24,61,120,170,193,198,199,200,201,201,202,202,202,203,203,203,203,202,202,200,196,193,194,197,198,198,197,195,194,193,194,198,203,203,194,183,184,192,193,177,144,118,113,119,130,137,131,125,131,138,137,128,122,126,135,137,129,121,120,128,135,130,119,119,131,141,142,142,146,143,130,115,117,138,150,138,122,131,150,148,130,125,141,146,129,122,141,155,138,116,123,141,124,81,52,39,28,21,20,20,21,24,25,25,29,36,36,26,14,10,11,16,24,32,45,65,92,116,128,128,129,142,156,160,154,148,147,145,143,147,157,164,165,159,158,158,157,157,160,165,167,165,166,173,181,188,184,172,157,136,118,107,93,83,90,106,115,114,107,109,125,143,159,178,188,177,159,152,155,159,161,158,147,142,147,152,158,166,168,162,152,138,127,130,139,143,143,145,151,160,163,157,141,122,114,126,148,168,179,178,162,148,149,155,155,151,144,126,108,101,101,100,99,95,94,95,95,100,110,111,105,106,109,
86,86,88,88,86,88,90,79,62,62,75,89,96,99,103,115,128,128,121,116,112,109,107,105,101,99,103,109,99,64,29,14,12,17,43,97,157,190,198,199,200,201,202,202,203,203,203,204,204,203,203,202,199,192,187,189,195,198,199,198,198,197,195,193,196,202,203,195,184,182,189,191,172,134,110,114,127,140,143,131,121,128,140,139,123,112,122,140,144,129,117,121,137,142,131,118,119,132,138,134,132,134,131,121,114,121,137,142,129,122,136,151,142,123,123,141,144,127,122,141,154,141,124,134,151,134,90,57,40,28,21,20,20,22,26,29,27,29,37,38,28,16,13,15,20,25,30,34,43,61,82,103,117,127,141,154,157,150,143,143,145,144,143,149,159,164,160,157,161,161,158,157,162,166,161,159,168,177,178,174,164,147,128,115,111,105,106,122,144,154,148,129,114,118,133,153,176,187,175,156,152,162,170,172,165,153,148,153,156,158,164,169,163,147,131,124,129,137,140,138,136,142,154,160,154,142,131,125,128,140,158,173,179,174,160,149,151,159,161,157,140,120,106,98,96,97,95,95,95,93,97,105,104,104,112,117,
74,74,75,74,70,74,82,77,66,70,84,93,97,99,103,115,123,121,119,121,120,120,119,113,105,99,100,107,107,79,40,17,13,15,33,82,145,186,198,200,201,202,202,203,203,204,204,204,204,204,203,202,198,190,184,187,194,198,199,198,199,199,197,194,196,201,202,197,189,185,188,186,165,133,119,125,134,142,140,126,118,125,136,134,120,112,121,134,138,134,128,127,131,135,135,131,126,123,121,120,118,113,110,113,121,130,132,124,118,127,143,146,128,115,127,145,142,123,121,140,152,140,127,138,154,136,92,58,41,28,21,20,20,23,28,31,30,32,42,44,31,19,18,19,20,23,27,29,33,38,48,63,83,102,120,134,142,143,139,137,141,146,146,147,154,161,160,159,164,167,161,157,159,163,161,159,165,168,168,169,167,153,136,128,127,125,125,139,157,163,155,137,119,115,129,153,175,179,164,148,148,160,170,172,166,157,156,158,150,145,153,165,159,141,129,132,138,141,142,137,128,129,143,152,151,150,148,140,133,136,151,164,171,175,169,154,147,151,157,158,146,127,109,97,97,102,100,98,101,99,98,102,105,112,122,127,
71,72,74,71,63,61,67,69,68,78,90,96,98,99,103,112,113,105,107,119,125,128,130,123,110,100,98,106,110,90,50,23,17,18,30,70,129,176,196,200,202,203,203,203,204,204,205,205,206,205,204,203,199,192,185,186,193,199,199,198,198,198,197,195,196,200,201,196,190,189,189,181,156,132,131,138,136,136,136,128,118,119,129,135,129,116,111,118,133,146,144,131,121,127,144,149,137,121,116,121,119,107,104,117,134,143,132,115,114,136,155,148,124,116,136,156,147,124,121,143,159,148,129,134,151,138,96,60,41,29,23,22,24,29,35,36,32,35,47,47,32,22,22,23,21,20,23,26,28,30,32,38,51,69,88,106,125,142,149,144,140,147,155,156,151,150,152,158,164,165,160,158,161,166,167,167,169,170,170,175,179,172,158,151,152,150,146,150,160,164,158,146,129,118,131,159,177,172,155,140,139,150,160,162,159,156,160,157,137,125,139,157,152,133,127,135,144,150,151,141,124,121,134,143,149,158,161,151,142,142,152,163,172,179,176,158,141,137,143,149,143,125,107,95,99,107,103,101,109,107,98,98,108,121,129,132,
91,93,91,78,57,45,47,57,69,84,93,97,99,100,103,110,105,92,97,115,122,123,124,120,110,101,97,102,107,91,54,27,20,21,27,53,106,162,193,201,202,203,204,204,205,205,206,206,206,206,204,202,201,195,188,186,191,197,200,199,196,194,194,194,194,197,198,192,187,188,189,177,150,132,137,140,132,129,133,129,119,118,130,140,134,115,104,112,132,145,141,127,120,128,144,148,137,125,124,132,132,122,119,128,138,140,127,113,119,142,155,146,127,123,140,156,147,126,123,144,161,150,127,127,145,139,100,63,43,33,29,30,37,46,52,49,38,37,47,46,31,23,26,28,23,20,22,25,26,28,30,33,36,44,57,73,94,120,140,143,137,140,153,156,145,133,136,149,158,155,150,153,163,168,167,165,166,169,169,173,178,176,168,163,165,165,161,161,166,169,164,152,136,122,129,154,171,169,157,142,136,142,151,151,146,147,155,152,129,115,131,149,143,125,122,134,148,160,163,149,129,123,131,137,145,158,162,154,147,144,149,166,180,185,178,160,141,131,130,137,136,123,109,101,104,109,105,106,114,109,95,95,113,130,135,134,
119,119,111,84,52,37,41,56,75,89,95,98,99,100,103,110,102,87,94,114,117,109,106,106,104,100,97,98,102,90,58,31,22,21,22,39,86,149,189,201,203,204,205,205,205,206,207,207,207,206,203,201,200,198,194,191,189,191,197,200,197,193,192,193,194,195,195,190,186,187,186,171,146,135,139,135,125,126,134,131,121,119,130,138,133,120,114,118,124,129,131,131,129,128,129,129,131,135,139,142,145,143,139,138,133,123,114,117,132,147,147,136,129,135,147,150,137,121,125,146,158,143,122,125,146,143,105,68,50,44,43,47,56,66,70,62,47,39,41,38,26,21,26,29,24,20,21,23,24,26,30,31,31,33,38,46,58,78,101,121,131,138,146,149,142,135,138,150,156,153,150,156,166,168,164,161,161,162,161,161,165,166,162,160,163,165,165,165,169,169,163,154,142,129,126,139,157,166,162,146,134,135,144,147,141,142,152,152,134,121,131,143,137,124,125,139,154,164,166,156,142,135,136,137,141,150,155,150,142,135,142,164,180,182,173,159,147,136,127,127,126,120,117,119,122,121,113,111,114,107,94,97,120,140,143,141,
129,125,109,76,46,38,48,66,83,93,97,98,99,100,103,109,102,87,95,114,113,100,94,96,98,98,97,97,100,93,66,37,22,19,19,30,72,134,181,200,204,205,205,206,206,207,207,208,208,207,204,202,201,201,200,195,189,187,192,197,199,196,194,194,195,195,193,189,187,189,185,160,135,132,137,129,121,128,140,137,122,117,126,136,139,136,130,122,117,125,139,145,138,125,116,119,133,147,148,144,145,147,145,141,130,115,111,127,149,157,145,131,134,150,159,149,128,114,125,150,159,140,118,125,148,145,108,72,56,53,52,56,63,69,70,64,52,40,34,29,22,19,24,28,25,21,21,23,24,27,29,30,31,32,35,37,40,48,64,88,116,137,147,147,145,149,157,162,161,157,158,164,169,168,165,165,166,166,163,161,163,164,162,160,160,163,165,166,167,165,159,153,151,144,130,127,143,162,165,151,133,127,138,149,148,149,158,161,150,135,132,136,134,131,138,151,159,160,157,152,146,142,140,138,133,133,137,136,131,125,132,153,168,168,160,150,147,146,135,123,116,115,121,133,142,140,123,108,101,95,90,99,124,145,151,149,
112,107,88,59,40,44,60,77,89,95,97,99,99,100,104,110,103,88,96,114,111,96,91,94,97,98,97,96,99,98,80,50,26,17,16,23,54,111,168,197,204,205,206,207,207,208,208,209,208,208,206,204,203,204,203,198,192,190,189,192,197,199,197,195,194,193,193,192,191,193,183,152,127,130,135,123,117,128,140,138,124,116,122,132,139,140,134,125,122,130,143,146,140,129,120,121,133,142,142,139,138,136,134,133,131,125,126,138,152,153,142,134,142,159,161,144,122,116,133,158,161,137,115,124,147,146,113,77,58,52,50,51,54,57,57,57,55,44,34,30,25,21,26,32,32,29,29,31,33,34,35,36,38,42,44,43,42,43,50,65,89,115,132,138,142,151,161,163,156,150,150,158,163,160,157,161,167,170,168,164,164,167,167,164,161,161,165,167,165,159,151,147,150,150,134,121,132,157,169,161,140,126,135,152,160,163,168,172,167,147,129,129,134,139,148,159,162,154,140,133,134,139,144,140,126,112,109,114,117,115,118,133,147,150,142,134,141,152,142,119,106,108,118,132,144,145,125,96,79,77,81,95,118,139,146,146,
81,77,63,47,42,55,73,85,92,95,98,99,99,100,104,111,105,91,98,114,109,94,90,94,98,99,98,96,97,101,95,68,35,17,14,18,40,93,156,195,205,206,207,207,208,209,209,209,209,208,207,206,206,206,205,202,200,197,192,190,195,200,199,193,189,190,194,195,194,191,174,142,127,137,138,122,114,122,133,137,131,120,115,119,128,134,135,132,127,122,125,133,141,140,130,120,119,125,134,141,139,132,127,126,131,141,146,145,140,133,130,137,152,161,152,131,117,126,151,169,159,130,112,127,153,156,129,94,70,60,58,61,65,64,62,65,67,59,51,50,44,35,39,51,57,58,57,57,57,55,53,57,63,68,71,71,66,64,67,71,79,96,114,128,139,150,157,156,149,140,139,149,156,153,149,153,163,170,169,165,164,166,168,169,166,165,168,170,165,156,148,143,147,149,135,118,122,148,169,168,148,132,138,157,170,173,175,180,177,153,131,132,142,150,154,159,160,148,128,114,118,135,149,144,121,98,91,101,111,107,102,110,122,125,118,119,138,155,145,118,101,101,110,120,132,139,123,89,66,68,79,92,109,123,126,125,
56,54,48,45,52,68,83,90,93,95,97,99,99,100,104,111,107,94,100,114,107,92,89,94,98,99,98,96,96,102,104,82,45,20,13,15,33,81,145,189,204,206,207,208,209,209,210,210,210,209,207,207,206,207,207,207,206,203,196,190,194,200,198,190,186,189,193,194,191,179,152,123,120,137,139,125,115,118,127,134,131,117,107,108,118,127,132,131,121,108,108,123,136,136,125,112,108,116,131,141,139,132,126,123,131,146,150,139,124,115,119,135,151,153,137,116,112,132,158,166,147,118,109,131,160,167,148,119,96,85,89,101,107,101,91,89,93,93,92,92,82,66,69,88,104,107,103,97,92,82,80,93,104,107,111,114,110,104,103,103,103,112,125,135,144,152,158,160,154,144,142,152,160,159,156,159,166,170,170,167,166,166,168,173,175,173,173,173,169,163,158,158,160,157,140,117,114,137,162,164,148,138,148,166,176,176,176,182,180,161,144,141,148,152,153,156,157,147,130,116,119,138,154,148,122,98,94,107,115,107,95,96,100,97,94,108,137,157,152,130,108,98,101,108,119,131,124,94,69,73,90,101,107,110,107,104,
64,61,55,56,66,80,89,92,94,95,97,99,100,100,104,111,107,96,101,113,104,88,87,93,98,99,98,96,95,100,105,91,55,25,14,14,26,64,124,177,201,207,208,208,209,210,210,211,211,210,208,206,205,205,207,208,208,205,199,194,196,199,195,187,186,189,190,189,183,164,130,105,109,127,136,130,118,114,120,126,125,118,113,111,112,114,119,124,121,114,113,116,117,115,111,112,117,124,129,129,124,120,119,123,133,141,136,122,114,117,126,137,143,135,117,105,113,136,154,152,131,108,107,134,163,169,155,133,114,108,120,138,145,133,115,108,117,131,138,137,121,100,96,118,143,152,145,134,119,103,105,127,142,141,141,142,137,131,130,130,131,136,142,143,144,147,155,160,155,145,142,150,159,161,161,161,162,162,162,163,163,163,163,168,171,170,169,170,169,168,169,173,175,169,150,126,115,130,152,155,142,141,157,176,184,181,176,179,178,167,153,143,138,138,145,154,157,151,144,137,134,143,152,148,128,110,110,119,121,109,95,88,84,79,81,100,130,153,158,147,123,101,92,95,107,123,124,100,77,84,106,116,114,111,106,102,
101,94,80,74,80,87,92,93,94,95,97,99,100,101,104,111,107,96,101,113,102,84,84,93,98,99,98,96,95,97,103,98,69,34,15,12,19,45,100,162,197,207,208,209,210,210,211,212,212,211,208,204,200,199,201,205,207,206,203,199,199,198,190,182,182,186,187,186,179,155,121,103,110,124,133,130,117,109,114,124,129,132,129,119,108,104,113,127,133,133,126,113,103,103,114,128,137,136,127,118,112,109,113,127,139,137,123,113,119,137,150,149,138,120,104,105,124,148,157,148,125,105,110,138,163,167,153,132,115,115,132,149,151,137,118,110,122,145,160,160,145,122,110,123,151,170,172,161,140,122,124,146,162,165,160,151,138,132,135,141,145,148,145,137,135,142,151,155,149,139,135,140,148,153,155,153,152,153,154,154,156,156,154,155,158,159,159,161,163,165,169,174,177,174,162,143,126,126,138,142,136,140,158,177,189,189,180,175,170,159,149,139,129,128,140,152,152,148,148,147,141,139,139,137,130,121,121,125,120,109,96,82,73,71,76,91,115,137,149,150,134,108,90,87,97,113,116,97,82,94,114,121,118,116,114,113,
129,119,100,88,88,92,94,94,94,96,97,99,100,101,104,111,107,96,101,112,100,82,82,92,97,98,97,96,95,95,102,104,82,44,18,12,14,33,82,148,192,206,208,209,210,211,212,212,213,212,210,204,198,195,196,199,202,204,202,200,200,199,191,178,173,178,183,184,175,148,117,108,113,118,123,125,120,116,120,127,132,135,136,131,122,117,122,130,134,136,133,123,115,119,129,137,138,132,126,125,124,121,124,132,136,130,123,125,140,159,165,153,130,109,102,116,142,162,164,147,123,108,116,139,159,163,151,129,111,112,130,147,149,138,122,112,117,138,160,167,158,139,120,119,139,165,179,176,159,139,133,144,162,176,178,165,148,139,139,144,153,159,154,142,138,145,153,157,155,148,142,142,145,149,153,154,154,155,155,154,155,155,152,153,157,158,155,151,151,154,160,167,173,174,169,157,136,122,123,129,134,143,156,170,184,188,180,171,159,144,137,135,133,135,146,150,143,134,132,132,130,127,123,123,121,116,117,121,115,105,94,78,68,69,72,81,97,115,131,142,137,118,98,86,89,100,99,86,81,96,111,114,112,114,119,121,
134,124,105,93,92,94,95,95,95,96,98,99,100,101,105,111,106,94,100,111,98,80,81,91,97,98,97,96,95,95,99,105,91,56,25,13,13,25,65,127,180,203,209,210,211,212,212,213,214,214,212,206,201,197,195,193,194,196,195,192,195,201,198,184,173,174,177,176,165,138,113,108,108,105,111,121,128,130,128,123,121,128,141,150,147,136,127,122,120,126,137,143,144,143,137,128,122,122,132,147,152,146,139,132,124,123,134,151,165,170,161,140,117,104,112,137,161,173,166,143,117,107,118,137,154,162,153,132,113,109,120,139,150,147,136,121,113,123,146,159,156,145,129,117,122,142,161,170,165,148,133,132,146,165,178,176,166,157,147,143,151,166,169,163,157,154,152,157,163,163,161,158,153,152,157,161,161,161,161,161,161,160,157,157,162,164,157,148,142,143,149,157,165,167,165,157,141,122,116,124,137,149,156,163,172,173,170,166,152,136,128,130,137,146,153,151,139,123,112,108,111,112,108,108,107,102,104,113,113,104,92,79,69,69,70,74,87,104,121,133,134,127,110,93,87,91,89,81,80,91,106,110,105,108,122,130,
123,116,102,92,91,94,95,95,95,97,98,99,100,101,104,111,106,93,98,110,97,78,80,91,97,98,97,96,95,94,96,103,99,70,34,15,12,19,46,103,165,200,209,211,212,213,213,213,213,214,213,210,207,205,201,195,192,192,187,182,189,200,201,192,181,175,170,163,148,125,111,111,108,105,112,121,125,127,126,122,120,129,145,154,147,129,115,109,111,121,137,148,150,140,123,111,111,121,140,156,156,145,132,121,115,124,144,161,168,158,140,120,105,103,123,149,167,170,156,130,107,100,110,129,147,156,150,132,115,106,108,125,145,152,146,129,111,109,122,136,141,142,136,122,114,117,130,148,160,157,144,135,133,142,157,167,171,170,160,147,146,158,169,175,176,169,160,156,159,162,167,171,166,162,163,163,158,159,166,171,172,169,162,155,157,163,163,156,149,143,141,142,146,148,149,149,141,126,117,122,138,151,157,161,161,158,160,162,153,137,125,124,133,142,146,144,136,121,104,91,91,96,97,99,100,94,96,110,116,110,99,86,75,72,70,70,83,103,115,118,120,121,112,97,94,102,104,94,86,90,103,107,100,105,127,139,
100,97,91,86,88,92,94,94,95,97,98,99,99,100,104,110,105,92,97,108,95,76,78,90,96,98,98,97,95,93,94,101,104,82,44,18,13,16,36,87,152,195,209,211,212,212,211,210,211,213,214,212,211,211,209,205,202,199,189,182,188,196,196,193,185,172,160,151,132,109,106,112,111,107,109,111,109,109,113,116,119,123,126,123,110,93,86,91,98,105,112,114,110,100,87,85,95,107,118,123,116,104,95,91,94,108,122,129,126,113,98,88,83,89,107,125,133,131,117,97,82,79,90,109,125,131,125,110,98,91,92,106,126,138,135,121,102,92,97,109,122,134,137,126,111,101,104,124,150,162,159,147,131,122,126,138,153,166,165,152,142,140,146,156,168,172,165,157,149,146,151,158,162,164,165,158,146,144,155,166,171,169,160,146,140,145,155,159,154,144,133,124,120,124,133,141,141,130,118,118,133,150,160,162,158,156,162,166,159,143,129,124,124,122,122,128,129,119,97,75,72,88,102,107,104,95,95,108,118,117,110,99,86,78,70,67,80,97,101,95,94,97,94,88,99,123,132,118,100,97,106,105,97,103,122,131,
70,71,72,76,81,85,87,89,92,95,98,99,99,100,103,109,105,92,96,107,94,74,76,88,96,98,98,97,95,93,93,98,103,86,49,22,16,18,31,71,133,184,207,212,212,211,207,205,207,211,213,213,213,213,213,212,212,209,201,194,195,192,186,183,179,165,153,145,124,98,94,98,94,89,89,90,89,88,89,91,92,89,82,74,65,56,55,61,66,67,66,62,58,53,49,52,60,67,69,67,61,55,52,52,57,66,71,72,67,59,53,51,52,56,65,73,75,73,66,56,51,53,62,75,85,87,81,72,67,67,71,80,93,100,99,91,79,70,71,81,95,108,113,107,95,85,84,98,120,137,140,132,115,100,94,99,114,132,140,132,121,111,105,110,125,138,140,135,126,118,114,116,123,133,138,132,119,112,116,125,133,136,132,120,108,106,116,126,127,120,111,102,96,100,115,128,134,128,116,114,129,152,164,165,163,165,172,173,163,151,140,130,115,98,94,104,114,106,80,57,61,90,114,115,105,98,99,107,112,111,110,108,101,90,75,69,79,90,90,80,73,73,74,77,96,126,140,129,111,106,113,115,107,105,110,112,
42,45,52,62,70,72,74,78,85,92,97,99,99,99,102,109,106,94,98,107,93,73,75,87,95,98,97,96,95,93,92,94,98,86,53,26,18,19,26,53,108,169,204,212,212,209,204,201,202,207,211,213,213,213,213,214,215,213,208,204,201,192,179,172,167,160,155,150,128,100,91,92,88,86,87,86,85,79,71,65,60,56,51,45,42,40,40,41,42,40,38,37,36,35,35,36,38,39,39,38,37,36,36,36,37,40,41,40,39,37,36,37,37,38,40,42,43,44,42,40,40,43,49,54,58,58,54,50,51,55,59,64,68,70,70,66,62,60,61,65,70,75,80,80,76,72,71,74,83,93,99,96,88,79,73,71,79,92,99,96,91,83,73,71,81,93,99,98,93,87,79,75,79,89,93,90,83,75,72,74,80,83,83,77,68,63,68,75,78,76,73,71,70,75,87,101,110,110,103,104,127,154,164,163,162,167,172,169,157,147,141,128,103,78,71,80,90,84,63,47,61,97,119,111,101,105,110,109,103,95,97,107,112,102,83,73,78,86,85,76,67,65,68,74,87,107,119,117,110,107,115,123,122,115,109,105,
29,30,36,48,56,58,62,68,78,88,96,99,99,99,101,109,112,107,109,112,95,75,76,86,94,97,97,95,94,93,91,92,95,87,59,31,19,17,20,38,89,155,199,211,211,208,204,199,198,202,207,209,209,209,210,211,211,210,206,203,203,196,181,165,156,156,160,157,140,121,118,121,121,122,123,119,109,93,77,63,53,50,48,43,41,42,42,42,42,42,41,42,43,43,43,43,43,43,43,44,45,45,45,44,44,44,45,45,45,45,45,45,45,45,45,46,47,49,49,49,49,52,55,57,58,58,55,54,57,61,64,65,66,66,65,64,65,67,68,68,65,63,67,71,72,71,70,67,66,70,75,76,75,73,68,66,69,75,77,77,75,72,65,60,65,73,76,76,75,72,65,61,63,67,68,65,61,56,51,51,52,52,51,49,46,45,48,53,54,51,49,55,61,68,80,92,98,95,89,98,131,160,166,159,152,151,154,149,136,126,116,100,79,65,62,65,68,67,57,50,66,99,116,105,100,115,122,115,98,80,80,97,109,103,83,69,68,74,78,73,66,63,65,70,76,85,94,101,105,104,107,116,121,122,121,119,
28,26,27,35,43,48,55,64,76,89,96,99,99,98,100,108,119,123,125,121,104,89,88,93,96,97,96,95,94,93,91,91,93,90,68,37,17,13,15,28,71,135,187,207,210,208,204,199,199,202,205,206,205,204,205,206,207,205,201,199,200,199,186,163,148,148,154,153,149,151,157,161,160,159,160,156,140,112,87,70,57,52,51,48,47,48,49,49,50,50,50,51,52,52,52,52,52,52,53,53,54,54,54,54,54,54,54,54,54,54,54,55,54,54,55,55,56,57,57,57,57,58,60,61,61,61,60,59,61,64,65,65,66,66,65,65,66,68,69,67,64,62,64,67,68,68,67,65,63,64,67,68,69,68,66,65,66,68,69,68,68,67,63,60,62,66,68,68,68,66,63,60,61,63,62,60,58,55,52,52,52,51,49,48,47,51,59,65,65,58,54,65,79,87,101,116,118,109,101,113,147,171,170,155,141,132,130,122,109,97,82,65,58,63,66,60,57,59,59,57,69,96,110,100,96,113,127,119,94,70,66,79,92,88,74,61,56,61,69,68,62,59,61,66,70,75,84,94,103,105,105,106,111,123,133,135,
31,26,21,25,31,38,48,62,79,91,97,98,98,98,99,105,115,123,125,121,113,110,110,108,104,100,97,95,94,93,91,90,92,91,74,41,17,10,11,20,50,108,170,203,209,207,205,203,205,207,208,207,205,203,204,204,203,199,195,191,192,195,188,167,146,140,142,143,153,170,178,176,171,167,167,169,152,116,86,68,56,49,47,48,49,51,52,53,53,53,54,55,55,56,56,56,56,56,56,57,57,58,58,57,57,57,57,57,57,57,57,57,57,58,58,58,58,58,58,58,58,58,59,59,59,59,59,59,60,61,61,61,61,61,61,61,61,62,62,61,60,60,61,61,61,61,61,61,60,60,61,61,61,62,61,61,61,61,61,61,61,61,60,59,59,60,61,61,61,61,60,59,59,59,59,58,57,57,56,56,56,55,54,53,54,59,69,75,73,64,61,80,102,109,120,136,140,133,129,139,161,173,164,147,131,121,111,97,85,80,71,55,52,65,70,61,55,58,60,60,70,88,96,87,83,98,116,113,87,64,58,64,70,72,68,60,55,58,64,64,60,63,70,73,72,73,79,88,97,104,107,105,106,117,128,131,
31,24,16,18,23,28,38,59,80,93,97,98,98,98,98,100,104,108,110,109,110,115,121,120,113,104,97,95,94,93,92,90,91,93,78,45,18,11,11,15,35,88,156,198,206,206,207,209,211,211,207,205,206,206,206,206,203,197,188,180,178,184,187,173,150,142,146,150,163,180,179,170,166,161,159,164,154,120,86,66,54,46,43,45,50,53,55,55,56,56,57,57,58,58,58,58,58,59,59,59,60,60,61,60,60,60,60,60,60,59,59,59,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,61,61,61,61,61,61,61,61,61,61,61,60,60,61,61,61,61,61,61,61,60,60,60,60,60,60,60,60,61,61,60,60,60,60,60,60,60,60,60,59,59,59,59,59,59,58,59,58,58,58,58,58,58,57,57,56,56,60,65,67,63,54,56,83,115,127,134,144,149,149,147,150,160,163,152,133,119,108,94,77,71,79,77,63,56,64,70,66,64,64,62,62,69,76,73,67,68,81,97,100,83,65,58,59,60,64,69,70,68,66,63,59,61,77,90,85,73,72,80,86,89,97,104,102,98,104,111,112,
25,20,12,14,18,22,34,57,81,94,97,98,98,98,98,97,97,97,97,98,100,105,111,116,112,103,97,95,94,93,91,90,91,95,85,56,32,24,23,25,41,88,151,191,200,203,208,213,214,210,205,203,206,210,210,208,205,200,189,175,167,172,182,177,159,154,163,170,179,186,175,163,161,158,155,162,158,133,101,76,58,46,40,44,51,56,58,59,59,59,60,61,61,61,62,62,62,62,62,62,63,64,64,64,63,63,63,63,63,63,63,63,63,63,64,63,63,63,63,63,63,63,63,63,63,63,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,63,63,63,64,64,64,64,64,64,64,64,64,63,63,63,62,62,62,62,62,61,61,61,61,61,61,61,60,60,59,59,58,59,59,56,49,42,49,79,117,142,153,158,158,157,151,147,153,159,150,128,106,92,79,68,70,80,79,66,57,59,64,68,70,69,64,67,73,70,58,54,62,73,85,92,85,69,60,62,64,65,72,80,83,78,68,63,70,89,100,86,70,76,91,93,88,93,100,95,88,96,106,108,
21,16,10,10,14,20,34,59,81,94,97,97,97,98,98,97,96,95,95,95,95,96,99,103,103,99,96,95,94,92,91,89,91,99,102,93,79,69,65,68,80,113,157,186,195,201,208,213,213,210,206,204,208,212,212,209,207,205,196,180,168,166,173,174,166,164,173,178,181,182,172,161,160,160,161,165,162,147,125,98,71,50,39,43,53,59,61,62,63,63,63,64,64,64,65,65,64,65,65,65,66,67,67,67,66,65,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,67,67,67,67,67,67,67,67,67,67,67,67,68,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,66,66,66,66,66,66,65,65,65,64,64,64,64,64,64,63,63,62,61,60,58,51,41,38,48,72,106,140,162,167,163,159,151,146,153,164,160,135,107,89,76,67,71,77,72,60,53,50,52,57,63,65,63,69,78,73,58,55,65,75,82,89,84,68,59,63,70,72,75,83,88,87,84,84,87,94,93,76,69,86,106,102,88,90,99,93,86,100,116,121,
19,15,9,8,10,17,34,58,80,93,97,97,97,97,98,97,97,96,96,96,96,95,96,96,97,96,95,94,93,92,90,89,91,104,126,145,148,137,129,133,141,156,174,187,194,202,208,211,212,211,206,203,208,212,212,208,205,203,198,187,173,164,166,172,172,169,170,168,166,169,166,159,162,166,166,166,162,156,145,125,95,62,42,44,55,62,65,66,67,67,67,66,66,67,67,67,67,67,67,68,68,70,70,69,68,68,68,68,68,68,68,69,69,69,69,69,69,69,69,69,69,69,69,70,70,70,70,69,70,70,70,70,70,70,70,70,71,71,71,70,70,71,71,71,71,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,69,69,69,69,69,69,69,68,68,68,68,68,68,67,67,66,66,65,65,63,60,50,39,39,51,69,93,121,148,161,161,158,156,155,160,167,163,144,121,103,87,73,74,75,64,51,45,42,42,47,54,57,59,65,74,73,64,64,75,80,81,82,76,63,55,58,67,73,74,78,86,95,107,115,111,98,82,70,75,100,116,104,84,83,93,91,89,103,120,126,
16,12,8,7,10,17,32,55,77,91,96,97,97,97,97,97,97,97,96,96,97,96,96,96,96,95,95,94,93,91,90,89,91,106,140,176,192,185,175,177,185,190,191,192,196,203,206,208,211,209,201,197,202,207,208,205,200,197,197,193,180,168,167,177,181,173,163,156,157,161,158,155,164,173,172,167,165,162,157,146,122,84,53,48,58,65,67,69,69,70,70,69,69,69,70,70,70,70,70,70,71,72,72,72,70,70,70,71,71,70,70,71,71,71,71,72,72,72,72,72,72,72,73,73,73,73,73,72,72,73,73,73,73,73,73,73,74,74,74,73,73,74,74,74,74,74,73,73,73,73,73,73,73,73,74,73,73,73,73,73,73,73,73,73,72,72,72,72,71,71,71,71,71,71,72,72,71,71,71,71,70,70,69,68,68,67,62,51,40,42,56,75,93,110,128,144,151,155,160,163,163,159,154,144,132,120,103,86,81,73,55,42,40,41,44,50,52,50,53,59,68,72,69,73,81,81,76,72,66,57,50,50,58,65,66,71,84,101,122,135,124,98,77,70,82,106,116,101,79,75,82,84,87,100,112,114,
10,8,6,7,9,16,30,50,71,86,94,96,97,97,97,97,97,96,96,96,96,96,96,96,96,95,94,93,92,91,89,88,90,106,139,175,195,195,187,187,194,198,197,195,198,202,205,207,207,202,193,191,195,200,202,201,197,194,196,196,188,176,173,182,187,176,161,158,163,162,149,146,161,174,174,171,168,164,161,157,142,108,69,55,61,68,70,71,72,72,72,72,72,72,72,72,72,72,72,72,72,73,74,73,73,72,72,73,73,73,73,73,73,74,74,74,74,74,75,75,75,75,75,76,76,76,75,75,75,75,75,75,75,75,75,75,76,76,76,76,76,76,76,77,76,76,76,76,76,75,75,75,75,75,76,76,76,75,75,75,76,76,76,75,75,75,75,74,73,73,73,73,73,74,74,74,75,74,74,74,73,73,72,72,71,70,65,53,42,46,61,84,105,116,123,133,142,147,153,159,158,149,139,134,130,124,111,96,82,64,45,36,38,43,47,52,51,46,46,52,63,71,73,75,80,78,71,64,55,47,44,48,53,56,55,62,80,101,118,125,113,90,74,71,81,99,107,97,79,72,73,74,80,94,102,102,
5,5,5,7,8,14,28,46,62,76,89,95,96,97,97,97,97,96,95,95,96,96,96,95,95,94,93,92,92,91,90,89,91,105,132,161,181,187,183,182,188,191,190,190,194,198,202,202,197,189,185,188,192,196,199,200,198,193,191,191,186,176,171,176,183,177,167,167,168,158,141,138,152,165,169,169,166,163,163,162,153,124,84,63,64,70,73,74,74,74,74,74,74,75,75,74,74,73,74,75,76,76,75,75,74,74,75,75,75,75,75,75,75,76,76,76,77,77,77,77,77,77,78,78,78,78,77,77,76,76,76,76,76,76,76,76,77,77,78,78,78,78,79,78,78,78,78,78,78,78,77,77,77,77,77,77,77,77,77,77,78,78,78,77,77,77,76,76,75,75,75,75,75,75,76,76,77,76,76,76,76,75,75,74,74,73,68,55,45,48,64,88,112,125,128,133,137,138,140,147,148,134,119,114,114,110,102,92,75,53,37,33,37,42,46,50,49,43,39,44,56,68,72,75,82,83,73,59,47,39,41,50,55,51,48,54,71,89,97,96,87,78,73,74,82,95,102,97,85,74,68,65,74,90,96,94,
3,3,4,6,7,15,30,44,52,64,81,92,95,96,97,97,96,95,95,95,95,95,95,95,94,94,93,92,91,91,90,89,91,104,129,152,169,177,178,177,181,182,179,180,185,187,187,185,179,174,179,188,192,195,201,204,201,189,179,175,173,169,167,170,175,174,168,163,155,143,135,139,152,161,163,164,164,165,165,165,158,132,93,68,67,72,75,76,76,77,77,76,77,76,77,77,78,78,81,86,88,85,81,79,78,77,77,77,78,77,77,77,77,78,78,78,79,79,79,79,79,79,79,80,79,79,79,78,78,77,78,79,80,79,79,80,80,81,80,80,80,80,80,80,80,80,80,80,80,80,79,78,78,77,77,77,78,79,79,79,79,80,80,79,78,79,80,79,79,79,79,77,76,76,77,78,78,78,78,78,78,77,77,77,76,75,70,58,47,50,65,88,111,126,132,137,138,135,132,135,133,115,97,96,95,85,80,81,72,51,35,31,34,38,44,51,52,45,40,42,53,66,73,82,96,97,79,59,47,42,43,50,53,48,44,49,61,73,74,68,65,67,70,74,85,101,108,101,86,75,69,65,75,93,96,92,
1,2,3,4,6,15,29,39,43,55,73,87,94,96,97,96,96,95,94,94,94,94,94,94,94,93,92,91,91,91,90,89,91,105,129,148,160,169,173,175,179,180,175,174,176,172,165,161,159,159,167,178,185,190,195,200,198,185,169,160,161,167,170,169,169,167,159,147,136,129,132,144,161,168,167,166,169,168,166,165,159,135,97,72,69,74,77,78,78,78,78,78,78,78,80,85,90,94,99,106,109,104,97,93,89,83,80,79,79,79,79,79,79,80,80,80,80,81,81,81,81,81,81,81,81,80,80,79,79,81,86,92,95,96,96,96,96,94,88,84,82,82,82,82,82,81,82,82,81,81,81,80,79,79,79,80,81,81,81,80,81,81,81,81,82,87,92,94,95,95,92,86,81,79,79,79,80,80,79,79,79,79,79,79,78,78,73,60,48,51,66,86,107,122,133,140,142,137,129,122,114,98,88,94,91,71,64,76,76,56,38,31,32,35,42,52,55,48,42,44,57,73,84,96,108,103,79,58,50,49,48,46,45,43,44,49,59,67,64,56,53,56,62,69,82,106,118,104,83,73,69,67,80,99,100,93,
1,1,2,2,5,12,23,31,41,57,73,88,98,99,97,95,95,94,94,94,94,94,94,93,93,93,92,91,90,90,90,89,91,105,128,146,155,163,170,174,179,180,174,169,165,159,151,147,147,148,149,154,162,170,178,183,185,180,166,154,154,163,166,160,156,155,146,133,125,125,131,143,162,171,167,167,171,169,165,164,159,137,100,74,71,76,80,82,81,80,80,80,79,80,86,99,111,116,117,120,121,118,115,113,107,96,86,82,81,81,81,81,81,81,81,82,82,82,82,82,82,82,82,83,82,82,81,81,84,92,103,112,115,114,114,115,117,114,106,96,88,84,84,84,83,83,83,84,83,83,82,82,83,86,87,89,89,86,83,82,82,82,83,86,94,103,112,116,117,117,113,103,94,87,82,81,81,81,81,81,80,80,80,80,80,79,74,61,49,52,67,86,105,119,130,140,145,141,128,112,96,85,88,100,96,73,64,74,74,56,39,33,33,36,45,53,52,45,40,45,60,80,95,104,106,94,72,56,55,57,52,46,44,44,45,50,63,74,70,59,53,53,58,65,78,104,120,108,88,74,65,67,87,105,100,92,
2,2,2,2,4,9,15,25,42,64,84,100,108,105,98,95,94,94,93,93,94,93,93,93,93,92,91,91,90,89,89,88,90,104,129,148,156,161,166,170,175,176,170,161,155,152,148,146,146,145,140,134,134,142,152,158,163,166,162,152,147,152,152,144,140,142,134,121,118,124,127,135,154,165,163,166,172,169,165,164,160,138,102,76,72,78,87,93,90,84,81,81,81,83,94,112,123,119,108,101,99,101,108,116,118,109,95,85,83,83,83,82,82,82,82,83,83,83,83,83,83,83,83,84,84,83,82,84,91,105,116,118,111,103,100,104,113,121,120,110,95,86,85,85,85,85,85,85,85,84,84,86,88,86,84,87,92,92,88,85,83,84,88,98,109,116,119,118,119,122,122,118,111,100,88,83,82,83,82,82,82,82,82,82,81,80,75,62,49,52,68,88,107,118,126,135,142,142,129,106,85,76,84,95,92,77,68,70,65,51,42,39,37,40,52,58,51,42,42,46,57,75,91,97,93,83,67,57,62,66,56,49,52,53,48,50,67,84,81,66,55,53,58,63,72,93,110,111,104,86,66,72,99,110,94,81,
2,2,1,2,6,10,14,22,42,70,94,111,113,104,96,93,93,93,93,93,93,93,93,93,92,93,93,93,92,91,89,88,90,104,131,153,160,160,162,165,168,169,164,155,150,151,150,150,150,149,143,132,123,123,130,134,137,144,150,146,140,141,143,139,138,139,128,114,116,123,124,130,151,165,168,174,176,171,167,166,161,140,104,78,73,81,98,113,110,95,84,82,81,85,98,116,117,96,72,59,56,60,71,88,104,110,101,89,85,85,84,84,83,83,83,83,83,84,84,84,84,84,84,85,85,84,84,86,96,107,106,92,74,61,58,64,78,95,109,110,98,87,85,86,86,86,87,87,86,85,86,90,87,70,56,60,78,93,92,87,84,86,94,105,108,100,92,87,87,93,100,107,114,109,94,85,83,84,84,83,83,83,83,83,83,81,76,62,49,52,69,91,112,122,125,130,140,143,130,104,82,73,76,83,80,71,65,64,56,47,45,45,41,43,56,64,54,46,48,50,50,60,77,84,82,75,62,57,69,73,59,51,58,59,51,53,69,86,84,67,52,52,58,61,66,80,93,102,110,96,73,78,101,101,78,65,
3,2,1,3,8,14,17,23,40,63,86,101,102,94,89,90,92,93,93,93,92,92,92,92,93,96,101,102,100,96,92,88,89,104,133,156,162,161,163,165,166,164,157,150,150,153,153,152,153,152,146,135,122,113,112,113,114,122,135,139,138,142,147,149,151,150,136,122,124,128,123,129,150,166,177,184,181,174,170,169,163,141,104,78,73,83,107,133,137,117,96,85,83,86,99,113,102,69,41,29,26,28,35,50,76,101,104,93,86,85,85,84,84,84,84,84,84,85,85,85,85,85,85,85,86,85,85,88,96,97,78,52,35,26,24,29,38,55,80,98,97,88,86,86,87,87,87,88,87,86,88,92,82,51,25,28,57,87,94,88,85,87,97,102,86,61,46,41,43,50,58,73,95,106,97,86,85,85,85,84,84,84,85,85,84,82,76,63,50,53,71,95,119,130,131,134,143,145,131,107,86,78,81,84,77,62,55,55,48,41,42,45,44,47,59,65,56,47,48,47,42,49,64,72,71,64,54,56,71,75,63,55,57,55,52,58,69,79,78,63,51,56,66,66,64,69,76,86,97,91,73,72,82,79,68,64,
2,2,1,3,9,15,18,23,33,44,58,75,84,84,84,88,91,93,93,92,92,92,92,91,93,102,114,118,115,108,97,89,89,103,131,154,161,162,165,167,166,162,152,146,150,154,152,150,149,148,143,134,120,108,103,102,103,113,126,138,146,150,151,153,157,157,147,137,137,131,120,126,144,160,174,183,179,173,172,172,165,141,104,78,74,85,111,145,159,143,117,96,86,87,99,110,94,56,30,22,20,20,21,28,57,93,105,95,87,85,85,85,85,85,85,85,85,86,86,86,86,86,86,86,86,86,86,88,95,87,56,27,15,13,14,15,18,29,58,88,95,89,86,87,87,87,88,88,87,87,89,93,79,42,12,14,46,82,94,89,85,87,95,93,65,31,15,13,18,24,29,45,75,97,96,87,85,86,86,85,85,85,86,86,85,83,78,64,51,54,71,96,123,138,140,144,149,145,129,110,95,87,91,95,86,63,47,43,38,33,34,39,45,51,61,66,56,44,41,38,35,40,51,59,60,54,49,54,68,76,74,67,58,50,53,65,75,82,79,65,56,66,78,76,64,60,67,78,85,79,63,56,59,69,85,94,
1,1,2,5,10,14,15,19,24,26,35,57,78,85,85,87,90,91,92,92,92,91,91,91,94,105,120,127,125,115,100,89,88,102,129,152,162,163,161,163,165,162,153,148,152,155,149,142,137,137,137,134,124,114,106,104,109,119,129,139,149,151,147,144,145,147,147,147,143,129,113,117,134,145,159,170,171,170,173,174,167,142,104,79,75,86,113,149,170,164,143,117,97,90,100,109,91,53,29,23,21,20,19,24,52,92,106,96,87,86,86,86,86,86,86,86,86,86,86,87,87,87,87,87,87,87,86,89,94,84,50,20,11,11,12,13,14,24,53,85,95,89,87,88,88,88,88,88,88,87,89,93,78,41,11,12,44,81,94,90,86,87,94,88,57,22,6,6,12,18,22,35,66,93,95,88,86,86,87,86,86,86,86,86,85,84,78,65,52,55,71,92,119,142,150,153,154,145,128,114,101,90,88,94,93,71,45,33,29,26,27,35,45,56,69,72,58,45,41,38,34,36,43,51,53,50,49,52,60,74,84,78,63,52,57,75,93,103,96,77,66,74,86,83,67,56,64,78,80,67,51,46,57,86,120,135,
1,2,5,10,14,13,11,14,18,20,31,59,84,91,87,84,85,89,91,92,92,91,91,91,94,104,113,114,112,107,97,88,88,101,129,155,166,163,157,159,164,163,157,153,155,155,148,138,131,128,130,134,134,126,115,111,118,126,128,132,139,140,137,131,126,128,135,141,137,118,103,110,123,129,139,156,166,170,173,173,167,144,107,81,76,87,114,150,172,174,163,141,116,99,102,108,89,51,27,21,20,20,18,23,52,92,107,97,88,86,86,86,86,86,86,86,86,86,87,87,87,88,87,87,87,87,87,89,94,83,50,20,11,12,13,14,16,26,54,85,94,89,87,89,89,89,89,89,88,87,90,94,79,41,10,12,44,81,94,90,86,88,94,88,56,21,6,6,12,17,21,34,64,92,96,88,86,87,87,87,87,87,87,86,85,84,79,65,52,55,69,84,112,146,163,164,160,149,136,121,102,83,74,81,88,72,44,28,25,25,29,38,52,68,85,84,64,49,48,46,41,41,45,51,54,51,49,47,52,71,87,86,76,69,72,87,108,120,112,90,74,75,82,81,68,57,61,70,68,54,45,51,76,113,146,158,
1,2,6,12,15,12,11,15,21,24,38,69,95,95,82,74,76,84,90,92,92,91,91,91,94,101,100,90,86,91,90,86,87,101,128,154,165,163,161,163,164,161,156,153,152,151,146,139,134,128,122,125,132,127,115,111,116,118,115,116,122,124,123,117,110,111,118,125,121,102,92,105,121,123,127,143,161,170,173,172,167,145,109,82,77,87,114,150,172,177,173,161,139,117,110,109,86,48,24,18,18,17,16,22,52,92,107,97,89,87,87,87,87,87,86,86,86,86,87,88,88,88,88,88,88,88,87,90,95,84,50,21,12,13,14,15,18,27,54,85,94,89,88,89,90,89,89,89,88,88,90,94,79,41,10,12,44,81,94,90,87,89,95,88,56,21,6,6,11,16,19,32,63,92,96,88,86,87,87,87,87,87,87,86,85,84,79,65,52,55,67,79,109,154,180,179,169,158,145,125,94,68,61,72,79,66,41,26,25,31,39,49,63,83,98,91,68,56,60,59,51,48,51,56,59,54,46,40,46,72,95,101,102,104,102,104,112,117,111,94,75,65,66,66,64,61,60,60,58,53,52,66,98,135,157,163,
2,3,6,10,13,13,18,29,36,35,47,78,101,94,74,62,65,76,85,90,92,91,91,91,94,98,91,74,71,81,86,85,87,101,124,145,154,159,165,169,165,157,151,148,147,144,140,138,136,128,114,110,116,114,106,103,105,104,100,103,107,109,108,102,98,102,113,121,115,96,85,98,118,124,122,131,150,165,171,172,167,145,108,82,77,87,114,150,173,178,177,172,159,140,126,115,87,47,23,17,16,16,14,21,52,92,107,97,89,87,88,88,87,87,87,87,87,87,88,88,88,89,89,89,88,88,88,90,95,84,50,21,13,14,14,15,17,26,53,85,94,89,88,89,90,89,89,89,89,88,91,94,79,41,10,12,44,81,95,91,88,90,96,88,56,20,5,6,12,16,19,31,61,90,96,89,86,87,87,87,87,87,87,86,85,84,79,65,52,55,67,77,110,162,193,192,180,167,152,123,82,53,54,69,76,63,40,25,26,39,52,60,71,89,98,87,69,64,72,72,61,53,54,62,67,59,44,35,45,79,112,121,127,138,138,128,118,107,100,90,71,54,50,52,56,61,62,64,73,77,74,83,114,145,158,158,
3,4,7,12,15,20,32,51,58,50,53,81,101,88,63,51,54,64,76,84,89,90,91,91,93,98,90,72,70,80,85,85,88,101,120,134,142,151,161,164,158,149,144,143,144,142,139,136,133,124,108,101,104,102,95,90,91,90,88,89,91,92,92,89,91,105,122,130,124,107,92,94,108,117,119,124,140,157,168,172,168,145,107,81,77,87,113,149,173,179,178,176,171,160,145,127,93,50,25,19,17,15,13,21,51,90,104,96,88,88,88,87,87,87,87,87,88,88,88,89,89,89,89,89,89,89,88,90,95,84,50,20,13,14,13,13,14,23,52,84,94,90,88,89,90,90,89,89,89,89,91,94,79,40,10,11,44,81,95,91,88,91,96,89,56,20,5,6,12,16,18,29,59,89,95,88,86,87,87,87,87,87,87,86,85,84,79,65,53,56,67,76,109,164,198,198,188,178,161,124,76,47,49,65,70,59,38,24,28,44,59,66,75,87,87,77,67,67,77,81,68,54,54,65,74,64,47,38,48,82,119,131,137,153,160,147,121,97,90,85,67,49,47,49,50,55,66,84,103,110,100,98,120,144,150,147,
5,6,11,17,22,28,43,66,73,58,56,80,95,78,50,39,43,52,63,73,81,87,90,90,93,97,90,74,72,82,86,85,89,101,115,125,135,146,150,147,141,135,134,138,141,143,139,134,131,124,110,103,104,102,93,83,77,75,73,74,77,82,85,87,96,112,125,128,124,116,106,99,99,105,112,121,136,154,167,172,168,145,107,81,78,87,113,149,173,179,178,177,176,172,163,143,103,56,31,23,19,15,13,20,51,89,102,94,88,88,88,87,87,87,88,88,88,89,89,89,89,89,90,90,89,89,89,90,95,84,49,20,12,13,12,11,12,21,51,84,95,90,89,89,90,90,90,89,89,89,91,94,78,40,10,12,44,81,95,91,89,91,97,89,56,20,5,5,11,15,16,26,56,87,95,88,86,87,87,87,87,87,87,86,85,84,79,65,53,56,66,74,104,159,195,198,193,188,172,132,80,48,46,54,55,46,33,28,33,47,63,75,83,86,77,66,60,60,69,76,67,52,49,63,77,72,55,46,50,76,109,127,138,156,163,143,108,83,79,78,62,48,47,49,47,53,76,103,121,126,115,105,116,135,142,141,
11,12,16,20,24,31,47,69,76,61,58,77,86,64,37,30,36,43,51,61,71,81,87,89,92,96,89,74,73,84,86,84,88,100,114,126,138,147,144,134,127,125,130,135,138,142,141,136,136,134,121,112,111,109,99,83,70,64,62,65,77,89,95,100,107,114,116,112,109,112,108,98,91,93,103,116,134,154,168,173,169,145,108,83,79,88,113,149,173,178,177,178,178,176,173,157,113,63,36,28,21,15,13,20,50,87,101,94,89,88,88,88,87,87,88,88,89,89,89,89,89,89,90,89,89,89,89,90,95,83,49,19,11,12,12,11,12,22,51,84,95,91,89,89,90,90,90,89,89,89,91,93,78,42,13,15,45,81,94,91,89,92,97,89,56,20,5,5,11,14,15,25,56,87,95,88,86,87,88,88,88,88,87,86,85,84,79,65,53,56,66,73,101,154,190,193,187,186,176,137,84,51,43,43,40,34,33,38,43,52,70,88,95,87,72,60,52,48,54,62,59,46,41,54,73,77,66,54,55,76,105,123,138,155,160,134,94,71,69,69,59,49,48,48,49,64,93,117,122,118,109,101,108,126,141,147,
18,18,19,20,24,34,51,70,76,63,59,74,77,52,28,25,33,39,44,54,65,77,85,88,91,96,89,74,75,86,87,84,88,103,125,144,156,157,151,142,134,130,133,139,143,149,150,146,146,142,131,124,123,118,106,86,70,65,66,72,89,103,109,113,116,112,105,100,99,102,98,86,82,89,98,110,130,154,168,173,168,146,110,84,80,89,115,149,173,178,178,178,178,177,177,165,120,66,37,29,22,15,13,21,50,86,100,94,89,89,89,88,88,88,88,88,88,89,89,89,89,90,90,89,89,89,88,90,94,83,48,18,11,12,12,12,13,23,51,84,95,91,89,90,90,90,90,89,89,89,90,92,81,53,30,30,53,82,93,90,89,92,98,89,56,20,5,6,11,13,15,27,60,90,95,89,87,88,88,89,89,88,88,87,86,85,79,66,53,56,66,74,104,158,190,184,168,165,163,131,83,52,41,38,35,31,37,49,55,57,72,94,100,88,72,60,50,41,41,48,49,41,36,45,63,76,72,61,62,84,110,126,138,156,163,138,99,75,68,66,61,56,52,49,53,76,109,126,119,103,91,92,106,126,144,151,
17,17,17,17,24,36,51,67,74,63,56,67,66,42,22,22,30,34,39,49,63,75,83,87,90,95,88,75,77,88,88,84,89,108,138,167,178,171,164,161,152,138,133,139,148,155,156,153,149,139,129,129,131,127,115,93,77,77,83,90,100,109,114,118,118,110,102,98,97,96,89,80,82,94,102,109,128,153,168,172,168,147,111,86,81,91,116,151,173,179,179,178,176,175,177,166,122,66,35,27,21,15,13,21,50,86,99,94,89,89,89,88,88,89,89,88,88,89,89,89,89,90,90,89,89,89,88,90,95,83,48,18,11,12,13,13,15,24,52,84,96,91,90,90,90,90,90,90,90,89,90,94,93,80,67,66,79,93,95,90,89,92,98,90,56,20,5,5,11,14,16,31,65,93,97,90,88,88,89,89,89,88,88,87,87,85,80,66,54,56,66,75,108,164,192,174,144,135,137,118,79,50,40,40,39,35,40,55,63,60,68,89,98,85,69,64,58,44,37,41,43,38,34,40,55,69,72,67,69,84,104,120,133,153,166,152,124,100,82,70,64,59,53,48,54,80,114,128,118,98,84,90,113,131,138,140,
12,12,11,13,21,31,43,58,66,58,49,52,50,32,17,17,23,27,35,48,64,77,84,86,90,94,88,75,79,90,89,84,89,109,139,168,178,171,165,166,159,138,125,128,139,148,150,149,144,129,119,123,127,128,120,100,84,87,99,105,106,108,115,123,120,109,102,101,101,98,90,84,89,98,102,110,131,154,168,172,168,147,111,86,82,92,118,152,174,179,179,177,175,174,177,167,122,65,33,24,20,16,14,22,50,86,99,93,90,89,89,89,89,89,89,89,89,89,89,89,90,90,90,90,89,89,88,91,95,83,48,18,11,12,13,13,14,23,52,85,97,92,91,91,91,91,91,91,90,90,92,98,107,110,108,108,111,109,99,91,90,93,98,90,56,20,5,6,11,14,17,33,68,96,98,90,88,89,89,89,89,88,88,87,87,86,80,67,54,57,67,79,115,171,196,171,135,119,120,109,77,48,40,44,44,42,49,62,67,63,68,87,92,76,63,66,67,52,41,41,41,35,32,40,57,70,72,71,72,77,88,101,114,135,157,161,151,133,104,76,62,53,46,42,50,77,111,129,127,110,94,98,119,131,127,123,
9,9,8,10,15,22,33,49,59,51,38,34,31,20,11,11,16,23,35,52,70,81,86,86,89,94,87,75,80,92,90,84,89,107,132,153,164,164,160,163,163,148,130,123,130,144,155,155,145,126,113,113,119,126,124,109,95,97,106,110,110,115,129,138,133,118,107,105,105,102,95,91,92,91,91,105,131,154,168,173,169,147,110,85,82,93,119,153,175,179,178,176,174,174,178,167,122,64,31,22,19,17,15,22,50,85,98,93,90,90,90,90,90,90,90,90,90,90,90,90,90,91,91,90,90,90,89,91,95,83,48,19,11,12,13,13,13,22,52,86,97,93,91,92,92,92,92,91,91,91,92,99,109,118,122,123,121,113,100,92,90,93,99,90,56,20,5,6,12,15,18,35,71,98,99,91,89,89,90,90,89,88,88,87,87,86,81,67,54,57,70,89,127,175,193,173,144,132,131,115,78,46,43,50,50,51,61,70,69,64,71,86,84,67,61,71,73,58,48,47,43,34,31,45,68,78,75,75,74,70,71,80,90,108,134,150,151,138,107,75,57,48,40,36,45,71,109,138,147,132,111,107,121,126,118,114,
10,9,8,8,11,16,28,47,56,45,27,20,16,11,6,7,13,24,41,62,77,84,86,86,89,93,87,75,81,93,90,84,89,107,130,149,165,172,170,171,178,175,156,137,139,161,177,174,157,133,115,110,116,128,133,125,115,112,113,116,122,134,151,158,149,130,113,103,97,95,95,96,94,84,78,92,122,151,168,174,170,147,110,85,82,93,119,154,175,179,177,175,173,175,179,168,122,63,29,20,18,18,17,23,51,85,98,93,91,91,90,90,90,90,90,90,90,91,90,90,91,91,91,91,91,91,90,92,96,83,49,20,13,14,14,14,13,22,52,86,97,93,91,92,92,93,92,92,92,92,93,96,101,106,109,110,109,104,97,92,91,94,99,90,55,20,6,7,12,16,19,38,74,100,100,91,89,90,90,90,89,89,88,88,87,86,81,67,54,57,73,100,138,172,182,170,157,155,155,130,83,50,48,56,55,53,62,70,66,60,66,76,69,57,65,82,80,65,57,54,48,37,34,52,78,86,81,83,79,63,56,65,75,88,110,128,129,115,91,70,60,53,42,36,41,66,106,143,157,145,123,112,116,117,113,112,
10,9,7,7,9,14,27,46,52,37,19,11,9,6,5,6,14,29,50,70,82,86,86,86,88,93,87,75,81,94,91,83,90,109,133,156,177,190,188,183,190,194,180,159,158,178,191,185,170,149,128,119,122,135,146,144,134,128,128,136,147,155,162,164,152,131,111,97,88,86,91,97,96,86,75,79,107,144,168,176,172,148,110,85,83,93,120,154,175,178,177,175,174,176,179,167,121,64,30,21,19,18,17,24,52,86,98,93,91,91,91,91,91,91,91,91,91,92,91,91,91,92,92,92,92,92,91,92,96,84,50,22,14,15,15,14,13,22,52,86,97,93,91,92,93,93,93,92,92,92,93,94,95,96,97,98,98,96,94,92,92,94,99,90,55,20,7,8,13,16,20,40,77,102,100,91,90,91,91,90,89,89,88,88,87,86,81,67,54,57,75,107,145,170,175,170,166,168,167,137,88,59,59,64,56,47,52,62,62,57,59,61,52,47,66,91,93,78,66,60,54,46,44,63,89,94,93,100,89,61,50,63,78,87,104,123,123,105,85,75,71,62,46,37,41,62,98,130,146,145,130,114,105,103,106,108,
10,9,7,6,7,12,25,41,42,27,13,7,6,4,5,8,18,35,58,77,85,86,86,85,88,92,86,75,81,94,90,83,90,109,133,158,182,195,192,183,185,191,186,172,168,179,188,186,180,166,149,139,139,150,162,157,142,136,145,161,170,164,155,150,143,126,105,92,86,83,84,88,92,90,77,71,94,136,167,177,172,148,110,85,82,94,120,154,174,178,177,176,175,177,180,166,119,64,33,23,19,18,17,25,55,90,100,94,91,91,91,91,91,92,92,92,93,93,93,92,92,92,92,92,92,92,91,93,97,85,51,23,15,15,14,12,11,21,52,86,98,94,92,93,93,93,93,93,92,93,93,93,94,94,94,95,95,95,94,93,92,95,100,91,56,21,8,9,13,16,21,42,79,103,100,91,90,91,91,90,89,89,88,88,87,86,81,68,55,57,77,113,155,181,186,183,180,179,171,135,88,67,71,70,55,42,43,55,62,59,59,57,48,46,66,94,104,94,77,65,64,66,70,88,106,104,105,114,100,66,56,76,97,107,121,141,141,116,95,90,86,69,47,37,40,57,82,107,129,143,137,116,98,94,98,100,
8,7,6,5,6,11,23,34,31,18,8,5,4,4,6,12,24,44,66,81,86,86,85,85,87,92,86,74,81,93,90,83,89,109,131,155,176,184,179,174,173,176,178,173,171,178,185,189,189,180,165,158,159,167,175,166,151,148,162,178,180,163,142,133,131,122,103,90,86,81,75,75,80,86,78,67,87,133,167,176,171,148,110,86,83,95,122,155,175,179,179,177,176,178,179,163,115,62,33,23,19,18,18,28,62,99,107,98,94,94,93,92,92,92,93,93,93,94,94,93,93,93,93,93,92,92,91,92,97,85,51,23,15,15,13,10,9,20,52,87,99,95,93,94,94,94,93,93,93,93,93,93,93,93,94,95,95,95,94,93,92,95,100,91,57,22,8,9,13,16,21,42,79,104,101,92,90,91,91,90,90,89,89,89,88,86,81,69,57,58,78,117,166,195,202,200,198,195,179,137,90,74,78,72,56,42,41,52,61,65,67,62,56,58,73,94,106,99,82,71,80,99,116,130,129,111,105,115,104,75,69,94,121,135,148,162,154,124,102,99,96,75,49,37,39,47,64,89,120,144,143,120,98,91,91,91,
5,5,5,6,7,13,25,32,25,12,5,3,3,4,7,15,30,51,71,83,86,86,85,84,87,91,85,74,81,93,89,82,89,111,137,161,176,178,176,174,169,165,168,170,172,178,185,194,197,188,176,171,174,179,182,175,168,169,176,182,175,154,133,123,121,116,103,92,87,81,71,65,69,78,77,70,90,135,167,176,170,147,110,86,84,97,124,157,176,181,180,179,176,177,177,158,109,58,30,21,18,19,19,32,72,112,120,111,108,106,102,99,97,96,95,95,95,94,94,94,94,94,94,93,92,92,91,93,98,86,52,23,15,15,13,10,9,20,52,87,99,96,94,95,95,95,94,94,94,94,94,94,94,94,94,95,96,95,94,93,93,95,101,92,58,23,9,10,14,17,22,43,81,106,104,94,92,93,93,93,92,91,91,91,90,88,83,74,64,63,78,116,162,191,198,197,197,195,180,142,101,86,85,75,59,45,42,50,60,72,76,67,62,66,77,91,100,95,81,74,90,125,153,163,146,112,95,101,97,79,77,104,135,154,165,169,152,119,97,94,93,76,53,42,41,43,54,82,116,139,141,122,102,92,86,84,
4,4,4,6,9,18,32,36,24,10,4,3,3,4,9,19,34,55,74,84,86,86,85,84,86,90,85,74,80,93,89,81,89,114,147,175,187,189,191,188,176,165,165,169,167,166,174,189,196,190,183,182,183,183,185,185,183,179,176,173,161,143,127,116,111,109,105,100,95,85,70,61,66,78,80,76,95,137,168,176,169,146,111,87,85,100,130,160,178,182,182,179,176,175,175,155,105,54,27,19,19,22,23,35,78,123,135,133,134,131,125,119,114,110,107,104,102,100,99,98,98,98,98,98,97,98,98,101,106,92,54,22,12,13,12,10,10,22,54,89,101,97,96,96,96,96,95,95,95,95,95,95,95,95,96,97,98,97,96,95,95,99,106,97,61,24,10,11,15,19,24,45,85,114,113,104,102,103,104,103,102,102,101,100,98,96,92,85,75,69,79,108,144,167,173,173,173,172,164,140,112,98,91,78,64,51,48,54,62,74,78,70,65,70,79,91,97,90,77,73,92,129,158,164,143,106,81,82,82,73,76,102,135,157,167,166,146,113,88,82,83,74,59,51,51,50,57,81,109,126,127,117,103,91,84,82,
4,4,4,5,10,20,34,38,25,10,4,4,5,6,13,26,43,62,77,85,86,85,84,83,85,90,84,73,80,92,88,80,89,115,150,176,188,196,200,194,179,169,169,167,153,138,143,165,177,177,176,178,175,173,180,189,185,171,159,152,146,133,116,100,95,98,100,99,94,84,70,61,71,88,87,78,96,138,168,176,170,147,111,87,87,105,135,165,179,183,182,180,177,177,176,154,102,50,24,18,22,26,28,39,81,127,145,151,159,160,154,149,143,137,133,128,123,119,117,115,114,114,114,115,115,116,118,121,125,107,61,21,9,10,12,11,12,25,59,95,107,103,102,102,102,102,101,101,101,101,101,100,100,101,102,103,104,105,105,105,106,112,120,110,68,27,10,11,17,21,27,49,94,128,129,122,124,127,128,127,126,125,124,123,120,117,114,107,92,78,80,103,132,151,156,156,156,156,153,139,116,99,87,79,73,66,64,66,66,70,78,80,80,86,94,101,99,85,72,76,98,127,146,146,124,89,66,64,64,61,68,93,123,146,157,157,139,110,86,79,83,81,68,60,59,57,60,78,96,104,109,109,101,90,84,83,
4,4,4,5,8,16,28,31,21,8,4,6,8,11,21,39,58,72,82,85,85,85,84,83,85,89,83,72,79,91,87,80,88,111,135,149,155,165,172,169,159,155,157,148,123,101,101,119,134,138,142,145,143,147,161,173,167,151,138,134,133,121,98,80,77,82,83,82,82,80,71,66,78,95,87,72,91,136,168,176,171,148,112,88,88,107,139,167,180,182,182,181,180,181,180,155,100,47,22,18,24,31,33,42,83,130,150,159,171,176,174,172,169,165,162,159,154,150,147,145,144,143,144,144,144,146,147,152,153,125,69,24,10,10,12,13,15,29,67,109,123,120,120,121,121,121,120,119,120,121,120,119,119,119,121,122,123,125,126,128,130,137,145,129,78,30,11,12,19,26,33,55,101,139,145,144,151,155,156,156,155,155,154,152,150,147,144,134,111,86,82,104,137,159,165,164,163,165,166,150,119,90,76,76,81,82,80,76,67,66,80,94,101,109,114,112,97,73,62,77,106,129,138,130,104,70,49,47,49,51,63,82,102,121,136,136,122,104,90,91,100,98,78,63,58,53,56,73,85,89,97,106,103,91,82,80,
4,4,4,4,7,13,20,22,14,6,4,9,15,22,34,52,70,80,84,85,85,84,83,83,84,88,82,71,78,91,87,80,87,102,109,104,102,108,121,127,123,119,118,105,79,61,60,69,77,83,90,96,106,122,139,143,134,127,124,125,125,112,86,65,61,65,67,67,71,76,75,69,75,84,75,63,87,136,169,177,174,152,115,90,89,107,138,167,180,183,183,183,183,187,188,161,102,48,25,23,31,40,42,53,93,141,159,162,173,181,182,182,181,180,180,179,177,174,173,172,171,171,171,170,170,171,172,177,175,140,76,29,14,14,17,19,22,36,79,129,148,145,146,149,151,150,149,149,150,151,150,149,149,149,151,152,153,154,155,157,159,165,170,145,85,31,12,13,21,31,39,59,105,146,157,160,169,174,175,175,175,174,174,172,171,170,167,155,125,92,84,108,147,175,183,180,179,185,189,168,122,84,72,74,81,85,84,75,62,62,81,100,111,118,120,108,84,59,51,71,104,127,131,119,90,57,38,36,41,48,58,69,78,91,106,108,99,93,95,105,117,111,87,67,57,48,52,72,89,95,102,108,105,92,80,76,
3,3,3,5,9,14,16,15,9,5,7,16,31,43,52,65,77,84,85,85,84,84,83,82,84,88,82,71,77,90,87,80,85,94,88,73,65,69,83,96,94,83,76,62,42,33,35,38,41,45,53,65,85,112,127,121,109,110,117,120,119,108,85,63,56,59,63,65,67,72,72,64,59,61,58,59,90,140,173,181,177,156,121,96,91,105,135,166,181,184,185,186,187,194,198,171,114,69,54,56,65,73,78,91,127,165,172,165,171,181,185,186,186,185,185,186,186,185,184,184,184,185,184,184,183,183,184,191,190,154,91,47,35,35,37,39,43,59,102,152,169,163,164,171,175,175,174,174,175,176,175,174,174,174,176,177,177,177,177,177,177,184,186,157,95,44,26,28,36,43,49,69,113,154,166,165,173,181,183,182,182,181,182,181,180,179,177,164,131,95,85,108,149,183,193,189,188,198,204,178,126,87,78,81,81,82,83,75,62,64,83,101,110,116,112,92,66,50,49,68,99,122,126,113,85,54,38,36,40,47,53,58,61,65,75,83,84,89,98,107,116,115,99,79,64,51,53,77,102,113,115,112,106,94,81,76,
2,2,3,6,10,14,13,10,7,6,12,28,49,63,70,75,81,84,84,84,84,83,82,82,83,88,84,75,79,90,87,80,84,90,81,63,53,55,67,79,75,60,47,35,24,22,26,30,32,37,46,61,82,109,124,118,107,106,111,114,112,104,88,70,60,60,64,66,68,70,66,55,48,47,51,66,102,148,175,180,173,155,128,106,97,106,134,165,181,185,185,186,188,196,201,183,144,116,112,118,126,132,137,149,173,191,183,166,169,181,186,186,186,186,186,186,187,187,186,186,187,188,188,188,188,187,189,197,200,175,128,95,86,85,87,89,92,106,139,172,178,169,172,182,187,187,187,187,188,188,188,188,187,188,188,189,188,188,186,184,184,190,195,172,125,88,78,80,84,87,90,105,140,172,175,165,171,182,185,184,184,185,185,185,184,183,181,169,136,99,84,99,135,173,191,190,191,201,205,179,130,96,90,92,87,85,89,84,69,69,87,101,108,113,105,80,56,49,56,74,100,122,128,116,91,66,51,44,44,47,51,56,54,49,56,72,83,91,97,102,108,116,111,92,71,54,54,78,104,116,115,112,109,101,87,81,
2,2,3,5,9,11,11,10,10,12,20,38,58,70,74,79,83,84,84,83,83,83,82,81,82,88,91,87,89,95,90,82,84,88,77,59,49,51,61,69,60,43,30,21,16,17,22,28,34,44,57,70,87,109,125,126,117,111,109,107,103,96,86,74,64,61,64,65,68,68,60,51,47,48,58,84,120,151,167,167,158,143,129,118,110,116,139,163,175,178,178,178,179,184,190,184,168,158,160,165,170,173,176,182,191,193,180,166,166,175,180,180,180,180,180,180,181,181,181,182,183,184,185,185,187,188,189,196,201,191,168,152,147,145,146,148,150,157,172,183,180,173,178,188,193,193,193,192,193,193,193,193,193,193,194,193,192,189,186,183,182,188,193,184,162,146,143,144,145,145,147,156,174,188,179,165,168,180,184,184,184,185,186,185,183,182,181,171,141,103,82,85,109,151,183,192,192,201,204,178,133,104,101,103,97,95,100,96,79,75,90,103,110,113,104,80,60,57,67,82,102,122,131,125,111,95,78,62,53,52,58,63,56,47,53,71,83,88,92,97,105,117,120,102,74,53,53,74,93,100,102,107,113,110,95,86,
3,3,4,6,8,11,14,18,23,28,35,48,62,68,72,77,82,84,84,83,83,82,82,80,80,87,96,99,101,101,93,83,84,84,71,51,41,44,58,66,53,33,20,14,11,13,17,24,35,52,71,85,98,114,126,128,121,114,109,104,95,84,73,65,59,61,68,69,66,64,59,52,47,50,69,103,133,147,152,149,136,122,119,124,126,131,144,156,162,163,163,163,163,164,167,168,165,164,166,168,171,172,173,175,176,174,167,160,160,165,167,168,167,167,167,168,168,169,169,170,170,171,173,175,177,179,180,183,186,185,179,174,172,171,171,172,173,176,179,180,176,174,179,186,189,190,188,187,187,186,186,186,187,187,189,189,186,182,178,175,173,175,177,176,171,169,169,171,170,169,170,175,182,183,172,160,162,170,173,174,175,176,176,174,171,169,169,162,136,101,82,83,99,139,182,197,194,200,205,180,135,108,106,105,97,97,107,105,88,83,95,106,109,107,101,91,79,75,82,92,101,112,118,122,128,127,109,88,74,72,80,84,76,66,66,72,76,78,86,97,107,121,128,109,77,54,51,66,81,86,91,102,112,109,95,86,
9,9,9,10,14,19,24,31,41,48,52,60,68,71,73,77,82,83,83,83,82,82,81,79,79,82,90,96,97,95,88,81,82,81,64,42,31,36,57,69,52,28,16,11,8,9,14,22,37,60,86,104,114,121,124,121,111,104,103,100,89,73,60,52,50,59,73,73,63,63,67,61,49,48,72,109,133,137,135,131,115,99,102,117,128,134,138,142,144,145,145,145,145,145,146,147,148,148,148,150,152,154,155,154,152,151,150,149,150,153,154,154,154,154,155,156,156,156,157,158,158,158,160,162,163,165,165,165,166,165,165,164,163,162,162,163,164,165,166,166,165,165,168,171,174,174,174,172,171,170,169,170,170,171,173,174,173,169,166,163,161,160,160,159,158,158,160,162,162,161,161,163,166,165,158,152,152,155,157,157,158,159,158,156,153,152,152,145,121,93,86,96,112,147,189,201,192,197,206,182,137,110,103,91,74,77,99,109,102,97,102,104,93,80,84,97,98,92,97,101,97,87,81,94,124,140,131,113,101,101,112,119,113,102,93,83,73,72,85,102,114,129,138,118,84,58,49,58,73,79,84,94,102,99,88,82,
28,28,26,24,25,30,35,43,52,56,58,63,67,71,75,79,82,83,83,82,82,81,80,79,77,77,78,79,80,80,78,77,80,78,58,35,24,31,56,72,52,24,13,9,7,8,14,24,39,64,95,119,128,126,119,108,94,84,85,87,81,69,56,47,45,56,70,68,58,66,79,73,55,47,63,93,116,121,118,111,96,80,82,98,111,116,118,120,121,122,123,123,123,124,124,124,125,126,126,128,132,135,135,132,128,127,128,130,133,137,140,139,138,140,142,143,143,144,145,148,149,149,150,151,152,152,152,152,151,150,150,150,150,150,150,150,150,151,151,152,153,153,154,156,157,158,158,157,156,155,155,155,155,156,157,159,158,157,156,154,152,152,151,149,148,149,150,151,151,151,150,150,150,149,147,145,144,143,143,142,142,143,142,140,140,141,141,133,109,87,90,107,122,152,192,202,191,196,204,181,136,109,94,68,42,46,78,107,113,109,109,98,70,46,56,86,101,99,104,110,95,63,45,64,106,135,136,123,112,114,130,145,146,136,123,106,86,78,92,109,120,136,147,128,91,60,45,51,67,75,78,84,91,92,87,84,
49,49,47,41,39,42,46,50,54,56,58,61,63,67,74,80,82,83,83,82,81,80,80,79,76,72,67,64,65,69,72,74,79,75,55,33,22,28,52,67,47,20,10,7,6,9,16,27,42,64,94,118,128,124,113,97,78,66,65,68,68,67,61,51,47,53,59,55,50,65,84,80,60,47,48,65,90,106,104,93,79,66,65,77,88,93,94,96,97,98,98,98,99,99,99,100,101,102,103,105,110,114,113,108,104,103,105,107,111,116,119,118,117,119,122,123,124,125,127,131,133,133,134,134,134,134,134,134,134,134,133,133,133,134,135,135,135,135,135,135,136,136,137,137,138,138,138,138,138,138,138,138,138,138,139,139,140,140,139,138,137,136,136,135,135,135,136,136,136,135,135,134,133,132,131,130,129,127,125,124,123,123,123,123,124,127,128,120,96,78,85,100,109,140,186,204,195,197,201,177,133,106,86,53,25,27,61,100,117,116,113,95,56,27,34,67,91,97,106,115,96,54,32,53,98,127,129,114,100,102,122,143,151,146,138,125,104,93,101,113,118,132,148,134,97,63,42,43,59,71,73,78,87,92,92,90,
53,55,55,53,54,57,58,58,60,62,64,64,65,69,75,81,82,83,83,82,81,80,79,78,74,67,57,52,56,65,70,73,78,74,54,32,22,27,44,53,36,15,7,6,7,10,17,30,45,63,86,106,115,112,102,87,71,61,57,55,56,63,65,58,51,49,48,45,44,60,81,79,60,44,36,46,77,108,109,91,73,59,55,65,76,81,82,83,84,85,85,85,86,86,87,87,88,88,89,91,94,96,95,92,90,89,90,92,94,97,99,99,99,100,102,103,103,104,105,107,109,110,110,110,110,110,110,110,110,110,110,109,110,111,111,111,111,111,111,112,113,112,112,112,112,112,112,112,112,113,113,113,113,113,113,113,114,114,113,112,112,111,111,111,111,112,112,112,112,111,111,110,109,109,108,108,107,105,104,102,101,101,101,102,104,107,111,102,79,64,72,81,86,122,179,205,198,198,202,177,132,102,79,46,20,21,51,92,114,118,114,92,52,23,27,55,83,95,108,116,96,54,34,58,103,127,121,100,81,83,104,124,133,137,137,128,111,101,106,111,110,120,139,136,106,70,42,39,54,68,73,77,86,95,94,92,
38,41,46,54,63,69,69,67,69,73,74,73,73,76,79,82,82,82,81,80,79,79,78,76,69,57,45,41,49,61,69,73,77,73,53,32,23,26,36,36,23,10,6,6,7,10,17,30,47,64,81,94,97,93,86,78,69,64,59,51,50,57,62,57,49,44,43,42,43,59,80,79,59,41,34,45,81,122,131,110,83,62,54,63,74,80,82,83,84,84,84,85,85,86,86,87,87,87,87,88,88,89,89,88,87,87,88,89,89,90,91,91,91,92,92,92,92,93,93,93,94,94,94,94,94,94,94,94,94,94,94,94,94,95,95,95,95,94,94,95,96,96,95,95,95,95,95,95,95,95,95,95,95,95,95,96,96,96,95,95,94,94,94,94,94,96,96,96,96,95,95,94,94,94,94,94,93,92,91,90,90,89,90,90,92,95,97,87,66,56,64,69,73,112,176,205,199,199,203,179,133,99,73,41,17,18,45,85,110,116,112,89,50,24,26,50,79,95,109,116,93,52,35,62,108,129,117,92,74,76,91,104,113,126,132,122,106,99,104,106,101,106,126,137,120,85,53,41,53,70,78,80,88,98,99,97,
21,23,31,45,60,68,69,70,74,79,81,80,80,81,82,81,80,78,74,71,72,75,75,70,60,44,33,34,45,57,66,71,76,71,52,31,22,25,30,25,13,6,5,5,6,9,16,30,47,63,77,87,87,79,72,68,64,60,55,50,49,53,54,49,43,39,40,41,43,58,80,81,62,45,39,50,87,132,150,136,106,75,59,64,76,81,83,85,86,86,87,87,88,89,90,90,90,89,90,90,90,90,89,89,89,89,90,90,90,91,92,93,93,93,93,92,92,92,92,91,91,91,91,91,91,91,91,91,91,91,91,91,91,91,92,92,92,91,91,92,92,92,92,92,92,92,92,91,92,92,92,92,92,92,92,93,93,93,92,92,91,91,91,91,92,93,94,94,93,93,93,92,92,92,92,92,91,90,90,90,89,89,88,89,90,92,92,80,63,58,67,69,72,111,174,204,198,198,203,179,133,97,69,36,13,13,40,80,107,115,110,85,48,23,25,49,77,96,110,113,89,48,34,64,108,126,113,89,74,74,82,91,103,119,124,110,94,90,97,99,94,95,117,140,136,105,70,48,52,71,82,82,87,101,108,108,
11,14,22,34,47,55,57,64,74,81,83,82,82,82,80,77,73,68,61,56,59,66,66,57,44,31,24,31,45,57,66,72,75,70,53,33,22,22,25,18,8,4,5,5,6,9,15,28,43,57,69,83,87,78,68,64,59,52,47,47,49,49,45,40,36,34,35,37,40,59,83,85,71,57,45,47,81,132,160,157,133,97,70,67,77,83,86,88,89,91,94,95,94,93,96,99,100,99,99,100,100,99,98,98,97,98,99,99,99,100,103,105,105,105,104,102,100,99,99,98,97,97,97,97,97,97,98,98,98,98,98,98,98,98,98,98,98,98,98,98,98,98,98,98,99,99,98,98,98,99,100,100,100,100,100,100,100,100,100,99,98,98,98,98,99,101,101,101,100,100,99,99,99,98,97,96,94,93,92,91,91,90,90,90,92,94,93,84,71,67,72,72,74,112,173,199,193,196,203,178,131,96,67,33,10,11,37,77,105,113,108,84,46,22,23,47,77,96,109,111,85,48,39,72,110,121,105,81,68,71,78,85,100,117,119,102,83,81,92,98,94,95,118,144,142,116,83,53,49,68,82,82,84,96,107,109,
10,13,20,28,36,39,44,57,73,81,81,79,77,75,71,67,61,53,43,39,44,50,49,40,29,20,19,31,49,64,71,74,74,66,51,33,20,18,18,13,6,4,6,7,7,8,13,22,33,44,59,81,92,83,71,66,58,46,40,42,44,41,36,32,30,29,30,31,37,62,89,91,78,66,47,39,71,126,162,168,154,118,82,71,78,85,93,99,100,103,110,114,109,103,105,115,122,124,124,125,125,124,122,122,122,123,124,123,123,125,129,132,132,131,128,126,124,123,122,121,120,120,120,120,120,120,120,121,121,121,120,119,119,120,121,121,121,121,120,120,120,120,120,120,121,121,121,121,121,122,124,124,124,123,122,123,123,123,123,122,121,120,120,120,121,123,123,122,122,121,120,120,119,117,114,110,105,101,99,98,97,97,96,97,101,107,111,106,92,79,76,72,73,111,171,196,190,196,204,179,130,94,66,33,10,11,37,77,104,112,107,83,45,21,21,46,76,97,108,108,84,49,47,84,119,120,95,67,56,64,76,84,96,114,117,99,78,76,89,99,98,103,126,146,137,114,87,56,45,59,75,81,87,94,97,97,
10,12,18,24,27,29,38,56,72,78,75,70,66,62,58,53,47,37,27,24,28,32,31,27,21,16,17,31,51,66,71,70,67,59,45,29,17,13,11,8,5,4,6,8,8,8,11,17,26,37,55,79,92,85,72,64,54,41,34,36,38,34,29,28,28,28,28,27,34,65,95,91,73,62,44,34,65,123,162,172,163,130,89,73,79,88,103,119,123,122,128,132,123,110,110,127,144,152,154,155,155,155,154,153,154,155,155,155,155,157,160,161,160,159,157,156,155,154,153,153,152,152,153,154,153,153,153,153,153,153,152,151,151,153,154,154,154,154,153,153,153,153,153,153,154,154,154,154,154,156,157,157,156,155,155,156,156,156,156,154,152,152,152,152,153,154,155,155,154,152,151,152,151,148,143,138,131,125,121,120,120,119,118,120,125,134,142,138,115,91,79,69,66,105,169,197,193,199,206,179,129,92,65,32,10,10,36,75,102,110,106,82,45,21,21,45,76,97,108,108,83,49,49,89,124,121,91,60,47,55,71,80,89,104,109,94,76,72,81,89,92,105,128,140,128,111,91,61,42,47,61,80,97,99,92,88,
9,10,13,17,20,25,40,62,77,79,70,61,55,51,45,40,33,24,16,14,15,17,18,20,19,14,16,28,44,54,56,57,57,53,41,24,12,8,6,5,4,4,6,7,9,12,17,22,32,47,63,78,87,82,68,55,45,36,31,34,38,33,27,25,27,30,30,26,32,64,95,87,62,48,34,31,65,124,164,174,165,133,90,73,79,90,112,138,149,145,139,133,122,107,105,124,149,166,171,173,173,173,173,173,173,175,175,175,175,177,178,178,175,174,173,174,174,174,174,174,174,175,176,176,174,174,174,174,174,174,173,173,173,174,175,175,175,175,175,175,175,174,174,174,175,175,175,175,176,177,178,178,177,176,177,177,178,178,176,174,172,172,173,173,174,175,177,177,176,175,174,175,175,172,169,165,160,155,153,153,152,151,151,153,157,163,168,159,129,97,80,67,62,101,166,196,194,200,206,178,128,92,66,36,16,17,41,77,101,109,105,83,49,27,27,49,78,97,107,107,83,47,43,82,120,121,94,64,47,48,61,73,84,97,101,91,77,69,69,73,83,100,120,129,126,118,99,66,41,38,52,78,100,100,92,90,
7,7,9,13,18,32,55,80,92,86,70,56,50,44,36,29,22,14,9,8,8,9,12,15,15,10,12,22,33,38,40,43,48,49,37,21,10,5,3,3,4,5,6,7,11,19,29,36,45,59,69,74,79,79,65,48,38,32,30,36,41,36,26,21,25,32,33,26,30,62,92,81,54,38,28,29,67,127,166,175,166,133,91,73,79,91,115,147,166,164,151,135,117,102,98,112,138,162,174,177,177,177,178,178,178,179,180,180,180,181,182,180,178,177,177,178,179,180,180,180,180,180,181,181,179,178,178,179,179,179,179,179,179,179,180,180,180,180,181,181,180,179,179,180,180,181,180,180,180,182,182,182,182,182,182,182,183,183,181,178,177,177,178,178,180,181,183,183,182,180,180,181,182,182,181,179,176,174,174,174,173,173,173,174,176,178,179,165,132,97,81,74,75,109,164,193,196,202,204,175,126,92,72,50,36,37,55,82,100,106,103,87,63,47,49,67,89,101,107,105,83,48,39,73,114,120,95,68,52,48,56,71,87,100,103,95,83,70,63,66,79,97,111,124,135,132,108,72,45,40,52,75,92,92,93,97,
6,6,8,14,27,51,80,103,109,95,71,52,43,36,28,20,14,9,7,6,6,7,11,13,11,7,9,20,30,33,32,34,38,39,32,20,12,7,3,4,6,7,8,10,15,27,42,50,54,60,62,62,66,68,57,42,33,27,29,37,42,36,24,18,22,32,34,26,29,59,85,75,50,36,27,31,72,130,167,176,167,134,91,74,79,91,115,149,171,174,167,150,130,111,101,105,127,154,171,176,177,177,178,178,178,179,179,179,178,179,180,179,178,177,177,178,180,181,181,180,179,180,181,180,179,178,179,179,179,179,179,179,179,180,180,179,178,180,181,180,180,179,179,180,180,181,181,180,181,181,181,181,182,182,182,181,183,183,180,177,176,177,178,179,180,181,183,182,181,179,180,181,182,183,183,182,180,178,178,179,179,178,178,179,180,180,179,165,130,96,84,88,101,127,160,182,191,197,194,163,115,82,70,60,54,55,65,78,88,91,91,84,73,70,78,94,106,108,106,101,82,53,44,75,115,119,91,62,49,50,60,74,89,99,100,94,83,70,64,66,77,91,105,126,144,141,115,80,54,48,60,79,89,89,95,100,
6,7,10,20,43,73,99,114,115,98,71,48,34,26,19,13,9,7,6,5,5,6,11,14,11,6,11,28,42,40,32,29,28,29,29,26,20,11,5,7,10,12,14,18,26,44,64,72,67,58,52,50,52,52,45,35,28,23,25,31,35,30,22,18,23,33,34,26,29,57,81,70,49,38,30,37,78,133,168,176,168,134,91,74,80,91,115,149,171,177,176,169,155,137,122,116,128,152,171,177,176,175,176,178,178,178,178,178,178,179,180,179,177,177,177,178,180,181,180,178,179,180,181,180,179,179,179,179,179,178,178,178,181,183,182,178,176,178,179,179,179,180,180,180,180,181,182,182,182,181,181,181,182,182,181,181,182,183,180,177,176,178,179,180,180,181,183,183,182,180,180,180,180,182,183,182,180,178,179,180,179,179,179,179,179,180,179,164,130,96,86,98,116,132,143,152,161,166,163,135,90,60,53,52,51,53,56,60,63,65,66,67,71,83,101,119,123,114,101,90,76,58,55,85,120,120,90,60,46,49,60,68,73,78,81,81,75,66,62,65,71,81,99,125,143,139,118,87,59,53,68,87,94,91,91,92,
6,7,11,26,55,86,103,107,105,90,65,41,25,16,11,9,7,6,5,5,4,5,9,12,10,10,21,48,65,54,34,25,24,26,30,31,26,16,9,11,17,24,32,42,54,72,95,102,87,66,53,49,48,43,36,31,27,23,22,25,27,27,25,24,32,43,43,33,37,64,85,73,54,45,38,44,82,133,167,177,168,134,91,74,80,91,115,148,171,178,179,178,172,162,150,142,145,159,175,179,172,165,168,175,178,178,178,178,179,180,180,179,177,177,178,180,181,180,179,178,178,180,181,180,179,179,179,179,179,177,176,177,184,191,187,174,168,173,178,179,179,180,181,180,180,182,183,183,182,181,181,181,181,181,180,180,182,183,180,177,176,178,180,180,179,181,185,190,189,184,179,178,179,181,182,182,181,180,180,181,180,179,179,179,179,180,179,164,130,96,87,97,113,122,121,119,120,121,119,101,67,42,37,39,40,41,43,44,45,46,47,53,73,103,131,147,142,117,91,73,63,58,64,95,124,121,95,68,50,45,51,52,47,49,61,71,70,63,60,63,66,72,88,113,130,132,119,92,63,54,67,86,95,91,84,82,
5,6,11,27,54,82,93,92,88,75,53,31,17,10,6,5,4,4,4,4,3,5,8,11,13,20,39,70,84,63,34,24,25,28,30,29,25,20,14,15,24,41,60,77,86,98,115,120,103,78,62,57,53,44,35,33,33,30,25,22,24,29,36,46,62,75,72,59,61,83,96,83,72,69,59,56,81,128,163,176,169,135,91,74,80,91,115,148,170,177,179,179,177,174,169,164,164,172,185,186,167,149,153,167,176,177,177,177,178,179,180,179,178,178,179,180,181,180,178,178,179,180,181,180,179,178,178,178,177,176,176,180,190,198,187,162,152,161,172,177,179,181,181,180,180,182,183,183,181,181,181,181,181,180,180,180,181,182,180,177,177,179,180,179,178,181,190,199,195,181,170,170,176,180,182,182,181,180,181,181,181,179,179,179,180,181,179,163,129,96,86,95,108,116,116,112,107,102,101,90,67,48,44,46,47,48,49,50,51,52,53,63,93,138,171,181,164,127,92,71,62,62,76,107,130,123,100,76,53,42,43,39,29,33,54,73,76,70,66,66,64,63,72,93,113,124,120,99,72,55,59,76,89,90,86,84,
5,6,10,21,43,66,77,77,72,59,38,21,11,6,3,2,2,3,3,3,4,6,11,17,23,36,57,77,80,59,33,24,27,30,27,23,23,23,19,19,30,53,78,94,101,108,116,117,103,82,69,64,59,46,36,35,39,39,32,25,25,34,52,76,103,117,111,99,100,114,113,99,100,107,97,79,84,116,151,170,168,135,91,74,80,91,115,148,170,177,178,177,176,176,176,177,180,188,198,194,166,139,142,162,175,178,177,176,177,179,180,180,179,179,180,180,180,179,179,179,180,180,180,179,178,177,177,178,178,180,183,189,199,200,179,147,134,144,159,171,178,181,182,181,181,182,183,182,181,180,181,181,180,180,179,179,180,181,179,176,176,179,180,180,178,182,195,203,191,166,152,157,171,179,181,182,181,180,180,181,181,179,178,180,181,181,178,162,127,95,86,98,116,129,135,137,133,126,122,117,102,90,87,89,89,89,90,91,92,93,95,103,130,168,195,200,179,141,112,97,88,88,105,131,142,130,103,74,52,46,50,41,25,28,54,80,90,84,75,70,65,58,62,81,102,117,120,109,86,62,56,70,86,92,92,91,
5,6,8,16,30,46,56,59,56,43,26,14,8,5,3,2,2,2,3,4,5,9,19,28,36,49,62,64,56,42,27,22,24,25,22,21,23,23,22,26,38,54,71,85,96,105,108,102,89,77,70,66,58,45,37,36,44,49,46,35,29,36,60,92,119,128,123,121,130,139,126,107,114,131,127,105,91,102,130,155,161,133,91,74,80,91,115,149,171,177,177,177,177,178,181,186,193,201,207,196,164,139,144,167,184,186,180,174,174,178,181,180,179,178,178,179,179,180,179,179,179,179,179,177,177,177,178,180,183,189,197,204,207,196,166,136,126,132,146,164,178,183,183,183,182,182,182,182,181,180,181,181,181,181,181,180,180,180,178,176,176,179,181,182,184,191,202,203,183,156,145,156,172,180,181,181,180,179,180,181,181,179,179,180,180,180,177,161,126,94,88,107,137,159,168,172,172,168,165,163,157,152,151,151,150,149,150,151,151,151,152,156,167,179,190,192,175,148,134,128,119,121,140,158,156,132,96,64,48,53,61,48,27,27,52,81,96,92,79,70,63,58,63,78,95,112,124,122,105,78,60,64,79,88,92,93,
4,5,7,12,22,33,43,49,47,34,20,13,10,7,4,3,2,3,5,7,9,16,32,46,52,56,55,43,33,27,20,16,16,17,19,22,24,23,26,36,46,50,58,72,87,96,94,83,71,65,65,61,52,43,41,42,52,65,67,54,38,36,53,80,97,99,97,105,122,133,119,98,101,118,122,107,90,90,109,134,147,127,89,74,80,92,116,150,172,178,177,178,181,184,185,188,193,196,190,170,139,123,139,170,191,193,178,164,165,174,179,180,179,178,177,178,179,180,180,179,178,178,178,177,176,177,180,185,191,199,203,203,196,174,142,121,117,123,136,158,177,183,182,182,182,182,182,182,181,180,180,181,181,180,178,177,178,179,177,175,177,181,185,189,193,199,202,193,170,149,149,168,184,187,183,179,178,178,179,181,181,180,179,179,180,179,176,160,126,94,90,118,159,186,195,197,198,197,197,196,195,194,193,190,187,186,187,188,187,186,186,186,181,171,165,164,155,139,133,130,124,127,144,159,154,125,85,53,43,52,59,44,27,30,48,75,93,90,76,68,63,61,64,70,84,108,129,135,125,98,68,56,63,75,84,88,
3,3,5,10,20,34,50,64,64,49,30,20,16,12,8,4,4,5,8,12,16,27,48,65,66,58,46,30,21,19,16,12,11,14,19,24,26,27,32,44,51,49,53,68,82,87,82,67,55,52,56,54,45,43,47,53,65,82,86,69,45,33,40,52,60,59,59,68,85,98,90,75,75,85,89,82,75,81,96,115,128,113,83,73,81,93,118,152,174,178,177,180,186,189,183,171,160,149,134,112,89,83,104,138,166,178,164,144,147,165,176,179,178,178,177,178,179,180,179,178,177,177,177,177,177,179,185,191,193,190,179,164,147,124,99,88,89,96,112,140,164,171,170,173,179,181,181,181,180,179,180,180,173,158,145,144,155,169,175,175,178,185,190,191,188,180,167,150,130,119,131,161,187,193,180,169,169,175,179,180,181,180,179,179,179,178,175,158,125,94,92,123,168,197,205,206,207,207,207,206,206,205,203,199,195,194,195,196,195,193,192,190,180,164,151,146,139,124,114,109,104,105,117,134,140,120,83,49,35,39,43,33,28,37,49,70,88,85,76,73,68,65,62,56,69,103,131,143,139,114,76,52,50,61,73,78,
2,3,4,10,21,39,64,86,91,73,48,30,24,20,13,8,7,8,12,17,23,35,56,71,69,56,39,22,15,15,13,10,10,16,21,26,29,32,37,45,49,49,54,68,78,79,70,53,41,41,46,46,42,43,50,61,75,87,87,69,45,31,28,31,33,34,35,41,54,63,60,54,56,60,57,52,57,74,89,101,107,95,74,70,81,94,120,153,174,177,177,181,189,191,174,141,106,80,65,55,48,50,62,83,117,147,145,126,129,154,173,178,178,177,177,177,179,180,179,178,178,177,177,176,177,181,190,193,179,152,121,96,78,63,53,50,50,55,72,105,136,147,147,157,170,175,177,179,180,179,180,179,158,116,84,84,113,149,166,171,179,188,188,176,153,126,101,85,74,70,83,118,158,177,164,147,151,167,177,179,180,180,179,179,178,178,175,157,123,93,92,124,169,199,206,207,207,207,207,207,206,206,204,201,198,197,197,197,197,196,195,193,187,177,167,158,143,124,112,109,107,106,113,128,138,126,89,49,27,26,26,24,33,46,54,72,88,84,82,85,78,70,61,48,59,97,131,147,144,117,77,49,44,53,61,64,
5,4,5,10,21,41,68,90,91,74,52,35,29,26,20,14,12,13,18,23,29,38,53,65,65,52,34,17,10,10,10,10,13,19,24,26,29,32,35,39,43,44,50,60,67,66,54,39,33,36,41,42,40,43,50,61,73,80,75,59,42,30,25,23,23,24,26,31,39,45,43,41,46,47,39,33,45,70,88,94,92,79,65,68,81,95,121,154,173,177,176,181,189,188,166,120,68,33,24,28,35,43,46,53,85,128,136,117,119,148,171,177,177,177,177,177,178,179,179,179,178,177,176,176,177,182,191,189,156,105,63,41,32,28,29,31,28,26,38,71,109,126,128,138,154,162,165,170,175,177,180,178,146,85,38,37,79,129,154,165,178,186,179,148,104,67,49,44,41,38,42,67,111,147,145,126,133,158,174,179,180,180,179,179,178,178,175,156,122,93,92,124,169,198,206,206,206,206,205,205,205,205,204,203,202,201,200,200,200,200,200,199,199,198,194,183,161,143,143,151,152,152,154,157,153,134,94,51,26,21,19,22,37,50,55,74,91,87,87,91,82,72,63,49,52,88,130,151,145,114,74,47,41,47,52,53,
10,9,7,10,21,42,68,81,69,51,43,38,35,33,29,24,20,21,27,32,37,43,51,59,60,51,33,15,7,7,10,12,15,20,23,26,27,29,30,32,35,37,41,46,50,46,36,29,32,37,40,40,39,41,47,55,63,67,61,49,38,31,26,23,22,22,25,29,36,41,38,36,39,37,28,24,39,68,88,91,84,70,60,67,81,94,119,150,170,175,176,180,185,183,160,114,57,20,14,22,34,45,50,54,84,129,140,120,120,148,170,177,176,177,177,176,177,178,178,179,179,177,176,176,178,183,190,183,140,77,34,20,18,19,23,26,24,18,25,57,98,120,120,125,135,141,146,155,164,172,178,176,141,74,24,23,67,119,146,160,176,182,168,127,71,35,29,38,41,37,31,41,82,128,135,117,123,152,173,179,180,180,180,179,178,178,175,156,121,92,92,124,169,197,204,205,205,205,204,204,204,203,203,202,201,201,201,201,200,200,200,201,203,206,205,196,177,165,175,189,194,194,194,185,165,137,99,61,39,34,31,32,44,51,53,73,92,88,85,88,80,72,66,51,48,79,128,155,147,114,74,47,40,44,48,50,
16,14,10,11,23,48,73,76,52,33,35,43,46,43,39,33,29,30,36,41,45,49,53,56,56,49,33,15,7,10,13,14,13,16,21,26,28,28,28,27,28,29,31,33,32,27,22,24,34,41,41,39,37,38,43,48,52,53,47,39,33,30,28,27,25,24,25,30,39,43,38,34,34,29,22,23,40,68,88,90,81,66,57,66,80,92,112,140,161,170,174,177,180,179,164,121,61,22,14,19,28,40,49,58,90,137,152,134,132,154,172,176,175,176,177,177,177,177,178,179,179,178,177,177,179,182,189,182,137,73,30,18,17,17,20,23,20,15,23,58,102,122,120,120,123,124,130,139,149,162,175,175,139,72,21,21,66,118,144,159,175,178,162,119,62,28,28,43,51,46,36,39,78,126,135,117,122,151,173,179,180,181,180,179,178,178,175,156,120,92,92,123,167,196,203,204,205,205,206,205,203,201,200,199,198,198,199,199,199,198,198,199,201,204,205,200,186,177,184,197,201,202,201,189,166,138,108,80,67,66,64,61,64,60,56,76,96,91,82,84,86,83,75,58,51,80,130,160,152,118,77,48,40,44,48,50,
25,21,14,12,23,49,75,76,48,27,31,46,55,54,48,43,40,40,43,45,45,46,46,46,45,39,27,14,9,15,17,14,10,12,19,26,27,26,25,25,24,22,23,24,20,15,14,22,35,43,41,38,36,37,43,47,46,41,35,31,29,28,28,27,26,25,27,33,40,40,34,30,30,24,20,27,48,75,89,89,80,64,56,66,80,90,104,124,141,153,164,172,177,182,177,137,72,28,17,20,24,31,40,53,90,143,164,152,149,162,173,176,176,177,178,177,177,178,179,180,179,178,177,177,178,181,189,186,145,79,35,23,21,19,20,22,19,17,27,62,106,125,122,120,117,114,119,127,138,155,172,176,139,70,19,19,64,117,144,158,173,178,166,125,67,30,30,44,52,48,37,42,83,132,139,121,126,153,173,179,180,180,180,179,178,178,175,156,120,91,91,122,166,195,203,204,206,208,209,208,205,201,198,197,197,197,197,196,196,196,197,198,199,201,203,201,193,186,188,193,195,193,189,179,162,140,118,102,97,98,97,92,86,76,73,92,113,104,85,84,97,103,94,71,58,84,134,164,158,128,90,58,45,47,54,57,
34,28,18,12,19,43,71,73,46,26,31,49,62,61,55,53,51,48,46,41,35,31,30,29,29,28,22,13,11,16,17,12,8,10,16,21,22,21,22,23,20,17,17,17,14,10,12,21,33,41,40,36,34,38,46,51,45,35,29,30,32,31,27,26,25,26,30,35,36,31,26,25,24,20,21,35,59,83,95,92,80,63,55,66,80,88,98,110,120,129,144,160,172,185,188,149,81,34,24,25,26,29,33,47,89,146,171,165,162,168,174,176,176,177,178,178,177,178,179,180,178,177,176,176,177,180,190,192,154,90,47,35,32,28,27,29,31,32,42,70,109,127,126,123,118,111,112,119,132,153,173,176,139,69,17,17,63,117,144,158,173,183,178,139,74,31,27,37,43,39,31,40,85,136,148,136,140,160,174,179,180,180,179,178,178,178,175,155,120,91,91,121,164,195,205,206,207,209,210,209,207,203,200,199,199,199,198,196,196,197,197,198,199,200,201,201,199,195,195,196,195,188,178,167,156,141,127,119,114,112,111,105,97,90,93,112,129,120,96,88,103,115,104,78,62,86,135,164,163,143,111,75,53,52,61,65,
33,28,17,10,13,34,62,67,43,26,35,57,71,68,62,58,54,46,38,29,20,16,16,20,25,29,25,16,12,14,12,8,6,8,11,13,14,16,18,18,15,12,11,10,8,7,10,18,29,36,36,33,33,37,46,52,46,35,30,37,44,41,34,31,30,30,32,33,29,22,18,20,21,20,27,44,64,86,99,96,82,63,55,65,80,88,97,105,108,111,122,140,159,179,186,150,82,35,25,28,30,31,33,45,88,146,173,169,166,171,175,176,177,177,178,177,177,179,179,179,177,176,175,175,176,179,190,194,159,99,62,53,49,42,37,41,51,59,64,81,111,129,131,130,124,116,114,120,135,157,175,176,138,68,16,16,63,117,144,157,173,187,188,148,77,29,21,29,33,30,25,36,83,139,160,157,160,170,177,179,180,180,178,177,177,177,174,155,119,90,90,119,161,193,205,206,207,208,208,208,207,205,203,202,202,203,201,199,199,200,201,201,201,201,202,202,202,201,201,201,198,191,179,168,159,149,140,135,128,119,116,114,109,107,112,123,133,129,112,101,110,119,106,84,73,94,135,162,167,156,128,87,57,53,59,62,
22,19,12,7,9,25,50,58,39,26,39,64,77,71,59,49,40,31,23,17,12,11,15,24,34,39,32,20,15,15,11,5,4,5,6,7,7,9,11,12,11,10,8,6,4,5,8,15,24,31,33,32,33,36,42,45,43,36,35,47,57,52,44,42,39,35,32,28,22,15,13,18,22,24,36,52,65,83,101,100,85,64,55,65,80,89,99,108,110,107,109,119,138,164,176,141,75,29,19,23,29,35,38,47,87,144,170,167,166,172,176,177,177,177,177,177,178,179,179,179,178,177,175,175,175,179,191,196,160,102,69,62,58,50,44,49,65,76,79,89,113,130,131,132,129,124,123,128,142,161,175,175,138,67,16,17,63,117,144,157,173,188,190,150,77,28,19,26,32,31,27,37,83,140,167,170,173,176,178,180,180,179,177,176,176,176,173,153,118,90,89,115,152,180,194,200,202,203,204,205,204,202,201,200,201,202,201,200,201,202,204,205,204,202,201,201,201,201,200,199,198,195,189,183,178,170,162,157,147,134,131,133,134,131,129,130,135,137,132,127,130,133,123,109,104,116,139,160,168,163,137,93,58,50,55,58,
15,13,10,6,7,17,39,49,35,26,39,61,68,58,42,29,21,15,12,11,10,12,19,31,41,42,32,20,19,19,13,5,3,3,3,4,4,5,5,7,9,10,8,6,5,7,11,17,23,29,31,33,35,37,37,36,36,34,38,55,66,58,47,44,41,35,29,24,19,13,11,16,20,25,39,53,61,78,98,101,88,68,57,65,79,88,100,113,117,112,106,105,116,142,159,130,67,23,14,19,28,39,43,51,86,141,167,163,163,171,176,177,177,176,176,176,178,179,179,179,178,176,174,174,175,180,192,194,157,97,62,54,51,45,41,46,60,71,75,88,115,130,127,125,127,128,130,135,144,159,173,175,138,68,17,18,64,117,144,157,173,188,190,150,79,32,24,30,38,42,39,46,87,142,168,171,175,178,179,180,180,178,176,176,175,175,172,152,117,90,89,111,138,156,166,174,181,185,188,189,187,183,181,181,183,186,187,187,188,191,194,197,196,194,192,193,195,196,194,192,192,194,195,196,194,190,186,182,172,160,157,159,158,151,142,137,136,138,143,146,146,148,146,142,139,139,145,153,157,153,136,100,64,54,64,71,
18,17,12,9,8,14,30,41,32,24,33,45,46,36,25,16,10,8,8,8,8,11,20,30,37,35,25,17,20,22,14,6,2,2,2,3,3,3,3,4,7,10,11,10,9,12,18,25,30,31,30,31,34,35,33,30,29,28,36,58,72,60,43,35,30,25,22,22,20,14,10,12,16,22,35,48,55,71,92,99,90,71,59,66,79,88,99,115,124,121,109,100,101,120,138,118,64,27,21,25,31,40,45,53,87,140,163,157,159,170,176,177,177,176,176,177,178,179,178,176,173,170,168,167,169,173,183,180,140,82,46,37,36,33,32,35,43,50,57,81,116,131,125,122,126,130,132,133,139,153,171,176,143,76,28,30,74,122,145,157,172,187,191,152,82,38,32,37,44,52,52,56,92,142,166,168,173,178,180,180,179,177,176,176,176,176,172,152,116,90,90,111,134,139,131,130,137,143,147,148,144,139,137,138,142,146,150,151,151,154,158,162,163,162,162,167,177,183,182,179,177,179,183,187,188,188,188,188,185,180,177,175,170,160,149,138,130,125,128,134,137,143,152,156,153,148,143,134,123,116,111,95,69,60,75,86,
29,25,17,12,10,13,25,35,29,20,22,29,30,27,22,17,11,7,5,4,6,10,17,24,27,24,17,14,19,22,15,6,2,2,2,2,3,2,2,4,8,14,18,16,13,15,22,29,33,32,29,27,27,28,28,27,26,26,36,61,77,61,38,28,24,21,21,24,23,17,12,13,16,21,31,41,49,66,85,93,88,71,59,66,79,87,95,110,123,124,113,100,96,107,123,108,64,35,33,34,35,39,44,52,88,140,161,153,157,170,176,177,176,176,177,177,178,178,176,170,161,153,150,150,150,153,159,154,117,66,34,25,24,24,24,26,28,31,41,73,115,132,127,127,129,130,129,129,136,153,173,181,156,103,66,70,104,136,148,156,172,187,191,153,85,42,35,39,47,56,57,61,94,141,162,165,171,178,179,179,178,177,177,177,177,177,172,151,115,89,89,115,144,141,109,90,91,96,97,96,93,90,90,92,96,102,106,107,107,107,109,113,115,114,116,126,141,150,150,146,142,141,145,149,151,152,154,157,161,164,166,165,162,155,146,135,121,109,105,109,116,127,141,151,150,142,128,105,78,65,67,67,57,54,70,82,
33,29,19,13,10,11,20,28,23,14,15,24,32,34,31,25,15,7,4,3,5,9,14,18,19,17,12,10,15,18,13,6,3,2,2,2,3,3,4,6,13,24,29,23,17,18,22,27,28,25,22,20,19,21,26,32,37,40,50,70,79,58,35,31,37,39,40,40,36,27,21,25,30,29,32,38,47,64,81,87,82,67,57,65,79,86,91,101,113,119,114,103,97,106,119,104,63,39,39,40,36,38,42,52,91,143,161,153,157,171,177,176,175,176,177,178,178,177,174,166,153,139,132,134,136,137,142,142,113,66,33,21,20,21,22,22,23,25,35,68,111,131,131,133,132,125,122,127,140,160,178,187,177,147,127,133,151,157,151,155,170,187,190,152,85,42,35,39,48,57,58,62,93,139,160,164,171,177,178,177,176,177,177,177,177,177,172,151,115,88,88,118,156,151,106,73,68,69,69,68,67,66,67,69,72,76,80,81,80,79,78,79,79,78,80,88,98,103,102,100,96,93,96,99,103,106,111,115,120,130,141,149,152,151,147,142,132,120,115,118,123,129,138,147,146,134,111,79,47,32,33,38,38,41,56,68,
28,24,16,11,8,8,12,17,15,10,14,27,39,41,35,27,17,8,4,3,4,7,11,14,15,12,8,7,9,11,9,6,4,3,3,3,4,6,8,12,20,31,36,29,22,21,24,26,25,19,14,13,13,16,27,44,56,61,69,78,72,50,35,42,57,65,66,65,57,47,46,56,58,49,44,44,49,64,79,83,77,62,54,64,78,85,88,93,100,107,108,103,100,110,122,106,64,38,38,40,37,36,39,54,97,149,164,154,158,172,177,176,175,176,178,179,178,176,174,168,156,139,128,132,139,139,145,152,127,76,37,23,22,23,23,23,24,28,38,70,111,130,131,133,130,120,118,128,145,164,179,190,191,180,173,177,181,168,149,149,167,187,191,152,84,41,33,38,47,56,57,60,92,138,160,165,172,176,176,175,176,177,178,178,177,177,173,151,115,88,88,120,162,164,118,78,68,73,77,78,78,76,75,74,74,74,76,77,77,75,74,73,72,71,72,75,77,77,77,76,75,74,75,79,86,98,109,115,120,131,146,159,167,169,170,170,167,163,161,162,162,158,156,160,157,140,108,69,37,22,22,26,27,32,48,60,
28,23,14,9,6,5,6,7,8,10,16,27,37,37,29,22,15,8,4,3,4,5,8,11,11,8,6,4,4,5,5,5,5,7,7,6,6,8,12,17,25,34,35,28,23,22,24,27,26,18,10,9,10,14,31,53,63,63,67,68,54,36,32,46,63,69,73,73,67,64,75,89,88,76,67,61,57,66,79,82,75,60,53,63,78,85,87,89,92,96,100,100,102,113,125,108,64,35,33,36,36,35,38,55,100,152,166,156,159,172,176,176,176,177,179,179,179,177,175,172,164,145,128,127,133,133,140,149,128,78,39,25,23,25,25,25,27,32,44,75,113,130,129,131,130,123,121,130,143,158,174,186,189,182,176,176,174,159,141,145,165,188,193,153,84,40,31,35,42,50,51,57,91,137,160,165,172,176,176,176,177,179,179,179,178,177,173,152,116,88,88,121,167,175,135,93,86,102,116,120,119,116,112,109,106,104,103,103,103,103,102,102,102,100,99,98,97,95,95,97,99,101,103,107,117,134,149,155,157,164,175,184,190,193,195,196,197,197,197,198,196,191,187,185,179,161,125,79,41,23,21,23,24,28,42,52,
44,36,20,10,6,4,3,3,5,9,16,23,29,27,20,15,11,7,5,5,5,6,7,8,7,5,4,2,2,3,4,4,6,10,11,9,8,10,14,20,29,36,34,24,18,17,18,21,22,15,8,7,9,14,31,50,52,46,48,49,35,22,23,36,49,54,60,63,60,63,81,97,98,91,88,80,68,70,80,83,75,60,53,63,78,85,87,87,89,91,93,96,101,114,126,107,63,34,30,33,33,35,38,52,95,148,165,156,160,172,176,177,177,178,179,179,179,178,176,173,166,146,120,107,105,106,114,124,109,69,37,25,24,26,27,27,29,35,49,79,114,130,129,131,134,131,129,131,137,151,169,179,178,170,163,160,158,151,144,150,169,190,195,155,86,40,31,34,39,46,47,55,90,136,158,164,171,176,177,178,179,180,180,179,178,178,173,152,116,88,88,122,169,182,149,113,115,142,163,169,168,166,163,160,157,155,154,154,153,153,152,152,152,149,144,139,134,132,132,135,141,148,153,157,164,175,184,186,185,188,194,197,198,201,203,204,204,205,206,207,208,207,205,203,198,183,149,96,48,24,19,21,22,24,33,39,
61,51,30,14,7,4,3,3,5,9,14,19,22,18,13,9,8,8,8,8,9,9,8,6,4,3,2,2,2,2,3,4,6,9,11,11,11,11,13,19,29,36,31,19,12,11,11,13,14,10,7,7,9,14,25,37,34,29,33,35,24,12,13,23,33,41,50,54,50,51,63,77,83,88,97,93,77,73,81,83,75,60,53,63,78,85,86,87,87,88,89,93,100,115,127,107,62,35,34,34,33,35,38,48,87,140,161,155,160,172,176,177,178,178,178,178,177,176,174,172,164,143,113,91,84,84,94,105,94,61,35,26,25,27,28,28,31,38,52,81,115,131,131,135,139,137,133,130,134,152,170,177,176,171,166,163,162,161,161,165,175,192,197,158,88,42,33,37,44,51,51,58,93,137,157,162,169,175,178,180,180,180,180,179,178,178,173,152,115,88,89,122,170,187,162,136,144,172,192,196,196,196,195,194,193,192,191,191,190,190,189,189,187,182,175,167,161,158,157,160,169,178,184,188,191,194,195,195,193,195,198,199,199,201,202,202,203,203,204,205,207,208,207,205,203,192,157,98,46,22,17,19,20,22,24,26,
71,60,36,16,7,4,3,3,5,9,13,16,16,12,8,7,9,11,12,13,14,14,10,6,4,3,2,2,2,2,3,3,5,8,10,12,12,11,10,15,23,28,23,14,8,7,7,8,8,8,8,9,10,12,17,21,20,19,24,24,15,7,8,14,23,37,50,54,48,43,43,50,60,77,97,99,82,76,82,84,76,61,53,63,78,84,85,86,86,86,87,90,99,117,130,109,63,38,39,39,34,35,38,46,81,132,154,151,158,171,175,176,177,177,176,177,177,174,173,170,161,139,109,87,79,80,92,104,92,60,35,26,26,28,29,29,32,40,55,83,116,131,130,132,134,132,127,124,133,156,174,179,179,179,177,176,176,175,174,174,178,192,198,159,89,43,35,41,51,59,58,62,95,138,158,162,169,176,179,181,181,179,179,178,178,178,173,151,114,88,89,121,169,188,166,145,155,177,189,192,194,196,200,201,201,200,200,200,200,200,200,199,198,194,189,183,179,177,176,178,183,189,193,195,196,196,195,194,194,196,197,198,198,200,201,202,201,198,195,193,194,194,193,191,189,179,141,82,36,19,16,18,20,20,19,19,
77,63,36,14,5,3,3,3,5,9,11,12,10,8,6,7,10,14,16,17,18,17,12,8,6,5,4,3,3,3,3,3,5,8,10,11,11,9,8,11,16,18,15,9,7,6,5,5,6,8,10,11,9,9,10,12,12,13,16,13,8,5,6,11,20,34,48,53,46,36,30,31,44,67,88,91,79,76,83,84,76,61,53,63,78,83,84,85,85,85,86,88,96,117,133,112,64,38,40,41,35,35,38,44,75,121,145,147,157,171,175,175,176,176,176,177,177,175,174,169,159,138,109,88,80,82,95,107,93,60,35,27,26,28,29,29,32,41,57,85,116,130,124,119,117,115,112,114,129,155,174,180,181,182,182,181,180,179,177,175,178,192,198,160,90,43,35,42,53,63,62,64,96,139,158,160,168,176,180,181,181,179,178,177,177,178,173,150,114,88,88,117,161,176,151,127,132,146,153,156,160,170,182,188,189,189,190,190,191,191,191,191,190,189,187,186,184,183,183,183,184,185,186,186,186,186,185,185,185,186,187,187,187,188,189,191,188,179,165,155,152,152,150,148,148,140,107,60,28,18,16,17,18,18,16,16,
82,67,35,12,4,2,2,3,5,7,9,8,7,5,5,6,9,14,18,20,20,19,15,12,11,11,10,7,6,5,4,4,5,8,10,10,8,7,7,9,12,13,10,7,6,5,5,4,5,9,12,11,8,7,7,7,7,8,8,7,5,5,9,15,23,31,40,43,38,28,20,20,31,49,63,66,67,74,83,84,75,61,53,63,77,83,84,84,85,85,85,86,92,113,133,114,66,38,40,40,35,34,37,42,69,111,136,142,154,169,174,174,175,176,176,177,177,176,175,172,164,144,113,89,79,82,97,109,95,60,35,27,26,28,29,30,33,43,59,84,114,127,119,109,104,101,100,105,121,148,170,179,182,183,182,181,180,179,177,175,178,193,200,162,90,43,34,41,53,63,62,64,96,139,155,156,165,176,180,181,181,179,178,177,178,178,173,149,113,87,86,112,150,158,124,93,89,95,99,102,108,123,140,149,151,151,151,152,152,153,154,154,154,153,153,152,152,151,151,151,150,150,150,151,150,150,150,149,149,149,149,150,149,149,150,150,147,134,114,98,92,91,90,90,92,88,69,43,25,19,18,18,18,18,17,16,
88,70,36,11,3,2,3,3,4,6,7,7,6,5,4,4,7,14,22,26,24,21,19,16,16,18,17,13,9,7,5,5,5,7,8,8,6,6,6,8,10,10,7,5,5,4,4,4,5,8,11,10,7,5,5,5,4,4,3,4,4,7,12,19,24,27,29,32,29,21,14,13,18,26,31,38,52,70,82,83,75,60,52,62,77,83,84,84,85,85,85,85,89,107,126,110,65,39,39,39,35,36,39,43,66,103,126,132,143,159,167,169,172,175,177,178,178,177,176,175,170,150,118,90,80,83,97,106,91,58,35,26,26,28,29,30,33,43,57,80,106,123,123,114,105,100,99,103,118,144,168,180,183,184,183,181,180,180,178,176,180,194,200,161,89,41,32,39,50,60,59,62,94,137,151,150,162,176,181,181,180,179,178,178,179,179,173,149,113,87,86,112,150,152,110,70,56,56,62,66,71,80,90,95,95,94,94,94,95,96,96,96,96,96,96,95,95,95,95,95,94,94,95,95,96,96,96,96,95,95,94,94,94,94,94,94,91,83,70,58,52,51,51,52,53,53,47,37,30,26,26,26,26,26,26,26,
87,69,35,13,5,3,3,3,4,6,7,7,6,5,4,4,7,15,26,33,31,26,23,19,19,21,21,17,12,10,7,5,5,6,7,6,5,5,5,7,8,7,5,4,4,3,3,4,5,7,8,8,6,5,4,3,2,2,2,3,4,7,12,17,21,22,22,22,21,16,11,9,10,12,13,20,40,66,81,82,74,60,52,62,76,83,84,85,85,85,85,85,87,99,112,98,61,39,39,39,37,40,46,50,64,93,112,117,127,143,154,158,165,172,177,179,178,178,177,176,171,152,119,91,81,89,103,105,85,54,33,26,25,27,28,29,33,41,54,71,94,117,128,123,113,107,107,109,124,150,172,181,183,184,183,182,181,180,179,178,181,192,193,154,85,40,31,37,46,55,55,59,90,132,146,146,160,175,180,181,180,179,179,179,179,179,174,150,113,87,88,117,157,156,108,61,41,41,52,59,59,60,61,61,58,56,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,58,58,58,58,57,56,57,57,58,58,57,56,54,51,46,44,42,41,40,40,41,40,39,38,37,38,38,39,39,40,40,
81,65,34,15,7,4,3,3,4,6,7,8,7,5,3,3,6,14,26,37,37,32,27,23,21,21,21,17,14,12,9,6,6,7,7,5,5,5,5,6,6,5,4,3,3,3,3,4,5,6,7,7,6,4,3,2,1,1,2,3,4,7,11,14,17,17,16,15,14,11,9,8,8,8,8,16,37,64,81,83,75,60,52,62,76,83,84,85,84,84,84,84,85,90,96,83,53,35,34,33,35,43,51,53,59,78,94,100,110,128,140,145,152,163,173,178,179,179,178,176,169,150,118,89,80,92,112,111,84,51,31,25,24,25,27,28,32,39,49,65,88,114,130,127,116,111,111,113,128,155,175,182,182,183,183,182,181,181,180,179,181,186,180,142,81,42,35,39,45,53,54,57,85,126,143,144,158,174,180,181,181,180,179,179,179,179,174,151,114,88,89,121,160,154,99,50,32,37,49,56,53,51,51,50,49,47,47,46,45,45,44,44,44,44,44,45,45,46,45,45,44,44,44,44,45,45,46,46,46,46,45,46,47,48,47,47,47,48,48,47,46,45,44,42,41,40,39,39,40,42,43,44,45,46,48,49,
80,64,35,17,9,4,3,3,4,5,7,8,7,5,3,3,5,11,25,39,42,37,34,30,25,21,19,15,13,12,10,8,7,8,7,6,5,5,5,6,6,5,3,3,3,3,3,4,5,5,6,6,6,4,3,2,1,2,3,4,5,8,11,14,15,15,13,12,11,9,8,7,7,7,9,19,42,69,85,86,77,61,52,62,76,82,84,84,84,84,84,83,83,85,88,76,49,30,28,29,34,44,51,51,54,70,83,88,99,117,130,134,139,150,164,174,179,180,178,171,158,136,106,80,69,81,102,104,78,46,29,24,23,24,25,27,31,36,47,66,94,119,129,123,112,108,107,110,124,151,173,181,181,182,183,183,182,181,180,179,181,182,172,134,81,47,42,45,50,56,56,59,85,124,140,142,158,174,180,181,181,180,180,179,179,179,175,151,113,88,90,121,153,137,79,35,24,31,42,45,42,39,41,45,46,47,47,47,46,46,44,42,41,41,42,43,44,44,44,44,43,43,43,43,43,43,43,43,43,43,44,45,46,46,46,45,46,48,49,48,47,47,46,46,45,43,41,40,40,40,41,40,41,43,46,47,
86,70,41,21,10,4,3,3,4,5,6,7,7,4,3,2,3,9,24,40,43,40,39,36,29,23,19,14,12,11,10,9,8,7,6,5,5,5,5,5,5,4,3,3,3,3,3,3,4,5,6,6,5,4,3,2,2,2,3,4,6,9,12,14,14,13,12,11,10,9,7,6,6,7,12,25,50,78,93,92,81,64,54,62,75,82,83,83,82,82,82,82,83,88,93,85,62,45,43,47,54,63,66,63,65,78,87,88,94,108,120,125,128,135,149,164,175,179,176,157,129,102,78,59,49,55,69,72,56,37,27,24,23,24,25,26,29,34,46,73,107,127,126,117,109,105,104,106,119,144,168,179,181,182,183,182,181,181,180,180,182,184,175,141,93,64,61,66,70,74,73,77,101,133,143,145,159,175,180,181,181,180,180,179,179,179,174,150,113,88,91,119,146,124,64,24,17,24,30,31,28,26,31,38,42,44,45,47,48,47,46,43,41,40,40,41,41,42,43,43,43,43,44,44,43,43,43,42,43,43,43,43,44,45,45,46,49,53,53,50,47,46,47,47,47,47,46,44,43,42,40,38,37,39,41,41,
92,78,50,27,13,5,3,3,4,5,6,6,5,4,3,2,3,7,19,32,36,36,38,35,30,24,19,14,11,10,9,9,7,6,5,5,5,4,4,4,4,3,2,2,2,2,2,2,3,4,5,6,5,5,4,3,2,3,4,5,6,8,11,13,13,12,11,10,9,8,7,6,7,10,15,29,56,86,102,101,88,68,56,62,75,81,82,81,81,81,81,82,87,98,107,104,91,81,82,86,92,98,97,91,92,101,104,98,93,98,107,114,118,122,130,146,162,173,170,140,94,59,43,35,30,31,35,37,32,27,25,25,25,26,26,27,29,35,48,78,115,132,127,119,112,107,105,107,119,142,166,179,182,183,183,182,181,181,181,182,187,194,191,168,133,113,111,116,120,122,123,128,144,163,165,160,165,175,179,180,180,180,180,179,179,179,173,148,112,89,91,120,149,129,68,23,13,16,18,18,17,17,23,30,35,37,41,45,46,47,46,45,43,42,40,39,39,40,41,42,42,44,45,44,44,43,43,43,43,43,42,42,43,43,44,49,61,72,69,58,53,54,56,57,57,58,58,58,57,56,54,52,50,50,50,50,
94,83,59,36,17,6,3,3,3,4,5,5,4,3,3,3,3,6,12,20,25,28,29,28,24,21,16,12,9,8,8,8,7,6,5,4,4,4,4,3,3,2,2,1,2,2,2,2,3,5,6,6,5,5,5,4,3,4,5,5,6,8,10,12,12,11,10,10,9,8,7,7,10,13,19,33,60,90,109,111,98,74,58,62,74,79,80,79,80,80,80,81,89,104,115,115,110,106,107,110,113,114,113,110,111,115,115,104,92,89,95,102,106,109,115,127,143,159,161,129,77,41,29,25,23,22,24,25,24,24,26,27,29,29,29,29,31,37,51,80,116,133,132,128,121,111,108,111,124,148,170,180,182,183,183,182,181,181,182,184,191,202,204,193,178,168,168,171,172,174,175,178,185,191,188,175,166,168,175,180,181,181,180,180,180,179,172,147,112,89,91,120,153,141,79,27,10,10,11,11,10,12,18,23,26,29,35,41,44,45,45,45,45,44,43,41,40,39,39,39,41,45,47,46,43,42,42,43,43,43,42,42,42,42,45,57,83,101,95,78,73,79,86,89,90,91,93,94,95,96,97,97,96,95,95,95,
99,89,67,45,23,8,3,2,3,4,4,4,3,3,3,2,2,4,7,11,14,17,18,18,17,15,12,9,7,7,7,7,6,5,4,4,4,4,3,3,2,2,1,1,2,2,2,2,3,5,7,6,5,6,6,5,5,5,6,7,8,9,10,11,11,11,10,9,8,8,9,12,15,18,22,36,63,94,113,118,106,81,60,61,73,79,80,79,79,79,78,80,86,97,104,105,102,101,102,103,103,104,104,104,105,107,106,98,88,84,87,91,95,99,104,113,127,142,146,126,90,61,46,37,33,32,35,39,38,32,28,28,30,31,30,30,32,38,51,80,116,135,135,133,123,112,108,113,128,154,174,181,182,182,183,183,182,182,181,184,190,195,193,186,180,177,177,177,177,177,178,180,181,182,177,163,149,152,168,179,181,181,180,180,180,179,171,146,110,88,89,114,147,141,85,31,10,7,7,7,8,10,14,17,19,21,29,38,43,44,44,45,45,45,45,44,44,42,40,38,40,48,53,49,43,41,42,43,43,43,43,43,43,43,46,66,99,120,113,97,93,103,113,119,122,125,128,131,134,138,141,144,146,147,148,149,
108,97,75,51,27,10,3,2,2,3,3,3,2,3,2,2,2,4,5,7,8,9,10,11,11,10,8,6,6,6,7,7,6,4,3,3,3,4,3,3,2,2,1,2,2,2,2,2,3,5,6,5,5,6,6,5,6,7,9,10,11,11,11,11,11,11,10,9,9,10,14,18,20,21,24,37,64,95,114,120,111,85,62,61,72,81,85,84,80,78,77,78,80,84,87,87,86,85,86,86,87,89,89,88,88,88,89,86,82,81,83,86,88,91,96,104,114,124,128,122,110,94,77,60,52,50,56,66,62,44,30,26,28,28,28,28,31,36,49,78,116,134,132,125,115,106,105,110,126,151,172,180,181,181,183,184,183,181,181,182,184,180,169,156,149,147,146,146,145,145,146,147,147,147,144,136,130,140,163,178,181,180,180,180,180,180,172,146,110,88,88,109,139,135,85,32,10,6,6,5,6,8,10,13,14,17,24,34,41,43,44,44,44,44,44,45,46,45,43,40,42,53,61,53,42,40,41,42,43,43,43,43,43,43,48,68,101,120,114,100,92,94,101,107,111,115,119,122,126,130,135,138,141,144,146,147,
116,104,79,53,29,12,4,2,2,2,2,2,2,3,3,3,3,4,7,8,7,6,5,6,7,6,5,5,5,6,7,7,6,4,3,3,4,4,3,3,2,2,2,2,2,2,2,2,3,4,4,4,4,5,6,6,7,9,10,12,13,12,11,11,11,11,10,10,11,16,21,23,24,23,25,36,60,90,111,118,110,86,63,60,71,82,89,90,84,79,76,76,76,77,77,77,77,77,77,78,80,81,81,80,78,78,79,79,79,80,81,83,84,86,90,96,103,108,109,109,109,103,88,74,66,64,73,86,80,53,31,24,25,26,26,26,29,34,47,77,116,133,126,116,107,101,102,108,121,144,167,179,181,182,183,184,183,182,181,181,180,174,162,149,141,138,137,136,136,136,136,137,138,138,137,134,135,146,165,178,180,180,180,180,180,180,173,148,112,89,90,114,144,135,82,32,13,8,6,5,5,6,8,11,13,15,20,28,36,40,42,43,43,43,43,44,45,46,45,42,45,58,66,56,41,37,39,41,42,42,42,42,42,42,47,67,97,114,111,94,75,66,67,70,73,76,78,80,81,83,86,88,90,91,93,94,
111,99,73,47,26,12,4,2,2,2,2,2,3,4,4,3,3,5,7,10,9,7,5,5,5,4,3,3,4,5,6,6,5,4,3,3,4,4,3,2,2,2,3,3,3,3,2,2,3,3,3,4,4,5,5,6,8,10,11,13,13,12,11,11,11,10,10,12,17,22,26,26,25,24,25,35,56,82,102,113,109,86,62,59,69,79,87,92,90,84,78,75,75,75,75,75,75,75,75,76,77,79,79,77,76,76,77,77,77,78,79,80,82,83,86,90,94,96,94,92,92,87,79,73,70,71,81,94,86,56,31,23,24,25,25,26,28,33,46,77,117,133,126,117,111,106,105,109,120,142,166,179,182,182,183,183,183,182,182,181,180,177,172,165,161,159,158,158,158,158,158,159,160,160,160,159,159,164,173,179,181,181,180,180,180,179,173,151,115,91,93,122,155,142,83,34,18,14,10,7,5,6,8,11,14,15,16,21,27,33,38,41,42,41,42,42,43,44,45,43,47,61,69,57,40,35,36,38,39,39,40,41,42,42,47,66,95,112,110,90,65,49,46,48,49,50,51,51,51,51,51,51,52,52,52,53,
86,77,56,37,23,13,5,2,2,2,3,3,4,4,4,4,3,4,6,9,9,7,6,6,6,5,3,3,3,4,5,5,4,4,4,4,3,3,2,2,3,3,3,4,3,3,3,2,2,2,3,4,4,4,5,7,10,12,13,13,12,11,10,10,11,11,13,18,24,28,28,27,25,24,25,35,53,75,91,102,103,84,62,58,67,76,83,90,94,90,82,76,74,74,74,74,74,74,74,74,75,76,76,75,75,75,75,76,76,77,77,78,80,81,83,86,89,89,86,81,76,69,65,65,68,74,89,101,88,57,31,23,23,24,25,25,27,32,45,77,117,135,132,130,127,119,114,116,127,150,171,181,182,181,182,183,183,182,182,182,181,180,180,178,177,176,176,176,177,177,178,178,179,179,179,179,178,177,179,181,181,181,181,180,180,179,175,154,119,93,94,126,162,148,86,38,23,20,16,12,9,8,8,11,15,16,15,15,18,23,31,37,40,40,40,41,43,44,44,44,49,64,73,60,42,35,35,35,36,37,38,40,41,42,46,65,93,112,110,89,62,45,42,42,43,44,44,44,44,44,44,44,44,44,44,44,
59,54,43,34,25,16,7,3,2,2,3,4,5,5,5,4,4,4,5,7,8,7,6,6,6,5,4,3,3,3,4,5,4,4,4,4,3,2,2,2,3,3,3,4,3,3,3,3,2,2,3,3,3,4,5,8,11,14,14,13,11,10,9,10,13,16,20,26,30,32,29,27,26,25,26,35,54,72,82,90,92,78,59,57,66,74,81,88,93,92,86,79,75,74,73,73,73,73,72,72,72,73,73,72,73,73,73,74,74,75,75,76,78,79,81,83,85,86,82,75,67,58,53,55,61,73,92,102,86,54,30,22,22,23,24,24,25,30,43,76,117,136,138,144,147,139,132,134,144,162,177,183,182,181,182,183,183,182,183,183,182,181,181,181,180,180,180,180,181,181,182,183,184,185,185,184,183,181,181,181,182,182,182,181,180,180,176,157,123,96,95,127,163,148,86,39,27,26,23,20,15,12,11,13,14,15,14,13,13,17,24,32,38,41,42,43,44,45,46,45,50,68,79,66,47,39,38,36,35,36,37,38,39,40,45,64,93,111,108,88,62,45,41,41,42,43,43,44,44,45,46,48,49,49,48,48,
55,52,46,39,30,19,9,4,2,2,3,5,6,6,6,5,5,5,6,6,7,6,6,5,5,4,4,3,2,3,4,4,5,5,5,4,3,2,2,2,2,3,3,3,3,3,3,3,3,3,2,2,2,3,5,8,11,14,14,12,10,9,9,12,17,23,28,31,33,32,29,26,25,25,27,38,58,74,80,80,78,66,53,54,64,73,81,88,93,92,87,81,77,74,73,72,72,71,70,70,69,69,69,70,70,71,71,71,72,72,73,73,75,77,79,81,83,83,80,73,63,53,47,49,54,65,83,93,80,51,29,21,22,24,24,24,25,29,42,75,116,137,141,152,163,162,158,159,165,174,181,183,183,181,181,182,182,182,182,183,183,183,182,181,179,178,178,179,179,180,181,182,184,185,185,185,183,181,180,181,182,183,183,183,181,181,178,161,127,97,94,126,161,146,84,39,28,29,28,26,23,19,17,15,14,14,14,12,12,15,21,30,41,51,54,49,46,45,47,47,53,72,84,71,51,44,43,41,39,38,37,37,38,39,44,63,92,110,107,87,62,46,42,42,42,43,44,44,45,46,48,51,53,53,52,51,
69,64,54,43,32,20,10,4,3,3,4,6,8,8,7,6,6,7,7,7,7,7,6,6,4,4,3,3,2,3,3,4,4,4,4,4,3,2,2,2,2,2,2,2,3,4,4,3,3,3,2,2,2,2,4,7,11,14,14,12,10,9,11,16,23,29,31,32,32,31,28,26,25,25,28,41,64,82,85,79,70,56,46,50,61,71,81,89,94,93,87,81,77,75,73,72,71,69,68,67,67,66,67,67,68,68,68,69,69,70,70,71,73,74,76,77,79,80,77,72,64,55,49,50,52,57,71,83,75,49,28,21,22,24,25,24,26,30,42,75,117,137,140,152,170,177,177,177,179,181,182,184,184,182,182,183,183,182,183,184,185,185,184,182,178,176,175,176,176,177,178,180,183,186,186,185,183,181,181,182,184,185,185,184,183,181,179,163,131,99,94,124,160,146,86,40,29,30,30,29,28,26,23,19,17,15,13,12,12,15,21,32,51,68,69,58,50,48,51,53,61,81,93,81,62,55,55,54,53,52,50,48,46,43,45,63,92,110,107,88,63,47,43,43,43,43,44,45,45,46,47,49,50,50,50,50,
78,72,59,46,33,21,9,4,4,5,6,8,10,10,9,7,7,8,9,9,9,9,9,8,6,4,4,3,3,3,3,3,3,3,3,3,2,2,3,3,3,3,2,2,3,4,4,3,3,3,2,2,1,2,5,10,15,19,18,14,11,11,16,23,29,32,32,31,31,30,28,26,25,25,29,44,69,89,93,84,69,52,41,46,58,68,79,89,95,95,89,81,76,74,73,73,71,69,67,66,65,64,65,65,66,66,66,66,67,67,68,69,70,71,72,72,74,75,74,71,66,58,53,53,54,55,64,76,71,48,27,21,22,24,24,24,26,31,43,76,118,137,140,153,173,184,186,186,185,185,185,186,186,185,186,186,186,186,187,188,189,189,190,186,179,172,172,173,174,175,176,178,184,189,189,186,184,183,183,184,186,187,188,187,185,184,181,166,134,100,93,122,159,148,88,42,30,31,31,31,31,31,29,25,21,18,14,12,13,18,29,46,70,87,85,72,65,66,72,80,90,107,118,110,97,93,93,94,95,94,93,90,83,69,59,68,93,110,108,89,65,50,47,47,46,46,46,47,47,46,47,48,50,52,54,55,
75,70,60,49,36,20,7,3,4,6,8,9,10,10,9,8,9,11,12,12,12,13,13,11,8,5,4,4,3,3,3,3,2,2,2,2,2,2,3,3,4,4,3,3,4,4,4,3,2,2,2,2,2,3,8,16,24,28,25,19,15,18,24,30,33,33,32,32,31,31,30,29,27,27,32,48,73,92,95,86,70,52,40,43,54,66,78,87,91,92,87,79,73,70,70,71,70,68,66,64,63,63,64,64,64,63,62,62,63,63,64,65,67,68,68,67,67,68,69,69,65,58,52,52,54,56,62,71,65,43,25,20,21,22,23,23,26,30,43,74,112,133,142,160,181,191,193,191,188,186,186,187,188,189,191,192,192,192,193,193,194,197,199,194,181,170,167,170,171,171,170,173,181,189,188,184,184,186,186,185,187,189,189,189,190,189,184,170,137,100,89,115,151,143,87,43,32,32,32,33,34,35,34,30,27,23,18,15,16,27,46,71,93,106,107,102,99,103,115,129,141,151,153,148,144,146,149,152,153,153,153,151,141,122,99,91,102,112,109,95,77,66,66,66,64,61,61,62,60,57,58,63,70,77,85,88,
56,54,51,47,36,18,6,4,6,9,11,12,11,10,10,10,10,12,13,13,16,18,16,13,9,7,5,4,4,3,3,2,1,1,1,1,2,2,2,3,3,4,4,4,4,3,3,2,1,1,2,2,3,5,12,24,33,36,32,25,23,28,34,36,35,34,34,33,33,34,37,38,38,37,41,56,77,87,85,78,70,55,41,41,50,61,73,79,79,79,76,72,67,65,65,66,67,66,63,60,58,59,60,61,61,59,58,57,57,57,58,59,61,62,62,61,59,60,62,64,61,53,47,48,54,59,63,65,55,36,22,18,19,20,20,21,24,30,42,68,100,123,144,169,186,191,191,187,180,176,177,180,182,186,190,192,193,195,196,195,195,201,206,196,175,159,154,156,156,155,154,156,163,171,168,163,167,177,182,183,185,186,185,186,190,190,184,169,138,100,86,106,133,123,78,43,34,35,35,36,38,38,37,35,32,29,26,23,27,45,73,98,113,125,139,146,145,148,161,176,185,187,182,176,176,181,186,187,188,187,183,179,178,170,151,130,120,117,113,107,102,100,102,103,101,98,98,97,91,86,89,98,110,123,134,139,
32,32,33,34,27,13,5,5,9,11,13,15,14,12,11,11,11,12,12,14,18,20,17,13,10,8,6,4,3,3,2,2,1,1,1,1,2,2,2,3,3,4,4,4,3,3,2,2,1,1,2,3,5,8,15,26,34,37,37,36,39,45,48,48,46,46,46,46,47,52,60,66,69,70,72,78,82,79,71,67,65,54,40,38,45,53,61,64,63,61,60,59,60,59,60,62,64,62,58,54,53,53,55,55,55,55,53,51,50,50,50,51,53,55,55,54,54,54,55,55,52,45,40,44,53,62,64,61,48,31,21,19,19,20,20,22,25,32,44,63,87,113,143,168,179,180,179,171,160,155,158,163,168,174,180,182,184,190,193,190,190,201,208,192,162,141,135,135,135,134,133,132,134,138,134,126,129,147,166,178,185,185,180,180,186,186,178,163,135,101,85,96,112,104,74,52,49,50,51,52,50,49,50,51,50,49,48,46,54,79,110,127,132,145,167,180,177,175,182,190,195,194,188,182,182,184,187,188,188,184,171,163,173,185,182,164,144,130,123,124,130,132,132,133,134,136,138,136,129,125,129,139,151,162,171,174,
26,24,19,17,13,6,4,7,10,12,15,18,17,14,12,13,15,16,17,20,22,21,17,13,11,8,5,3,3,3,2,2,1,1,1,1,2,2,2,3,4,4,4,3,3,2,2,1,1,2,3,5,8,12,19,28,35,41,50,64,77,84,86,87,86,86,85,85,86,93,104,113,119,120,118,108,89,71,62,59,58,49,36,35,40,45,49,52,51,49,49,50,52,54,55,59,63,62,58,55,55,55,53,50,49,49,48,48,46,45,44,45,47,48,48,49,50,51,52,51,46,40,37,40,49,58,63,59,45,31,25,25,27,30,34,37,41,47,57,71,90,116,144,163,170,172,170,158,142,136,140,148,155,162,168,170,174,182,186,183,187,202,211,195,161,138,132,132,132,132,131,126,124,124,118,102,95,110,140,169,188,192,186,185,188,187,177,162,137,106,89,94,109,113,102,94,95,96,98,96,86,78,85,95,99,99,99,99,107,129,152,158,151,155,170,177,171,161,157,160,165,165,160,155,153,155,160,167,174,172,154,142,157,181,188,181,166,151,143,145,150,149,146,147,152,159,164,164,161,159,162,169,175,179,183,184,
39,31,16,6,3,3,5,9,12,12,14,18,20,19,21,25,28,31,35,38,38,34,29,25,21,14,8,4,3,3,2,2,1,1,1,2,2,2,2,3,4,4,4,3,3,2,2,2,1,2,5,10,14,21,35,52,64,73,89,111,130,139,142,143,143,141,140,139,141,146,154,159,159,157,149,126,93,68,59,57,54,44,34,33,37,40,44,47,46,45,45,46,47,48,51,55,62,66,64,62,65,65,58,50,45,44,46,48,48,47,45,44,46,47,46,47,50,55,60,60,53,44,39,40,46,54,61,61,51,41,40,44,49,60,71,79,81,84,91,103,120,141,156,163,169,175,172,160,146,140,142,150,160,167,171,175,179,185,188,188,194,208,217,202,173,154,150,151,152,154,152,146,142,141,133,110,90,93,121,161,193,205,205,204,203,201,195,182,161,135,117,119,138,154,158,158,160,161,163,157,134,118,133,157,166,166,165,165,169,180,187,180,164,153,146,140,133,122,111,112,120,125,123,115,110,114,126,144,163,170,154,142,158,183,192,189,183,173,165,162,163,163,162,164,169,175,180,182,182,182,182,182,181,181,182,183,
45,34,15,4,1,3,8,15,18,18,20,25,30,37,47,55,56,62,73,81,81,77,73,68,59,43,23,10,5,4,3,2,1,1,2,2,3,3,2,3,3,4,4,3,3,3,2,2,1,3,7,13,20,35,62,92,113,126,139,154,166,173,176,178,177,175,175,177,179,183,187,185,178,171,160,134,100,76,69,68,64,52,41,38,41,44,47,48,48,47,47,47,48,50,52,54,61,67,67,67,70,72,65,55,47,46,49,52,55,57,57,56,60,63,62,60,65,75,86,87,76,60,50,51,60,68,73,75,72,71,77,84,91,105,122,132,135,137,142,152,167,178,175,167,173,182,182,175,171,170,172,177,184,190,195,198,201,203,204,205,209,217,219,205,185,174,173,175,177,180,180,177,173,172,164,144,123,118,134,168,201,217,221,222,221,219,217,211,199,183,165,158,171,191,200,202,203,204,206,196,166,145,165,195,205,203,200,200,203,206,201,186,168,149,127,111,108,104,95,97,111,124,127,118,110,113,126,146,167,176,162,150,166,190,197,195,191,185,175,164,164,171,177,180,183,188,191,192,192,192,190,186,181,179,180,181,
38,30,14,4,2,3,10,20,31,41,49,51,52,59,75,85,88,101,122,135,137,136,133,130,120,94,55,24,10,6,4,2,2,2,2,3,3,3,3,3,4,4,4,4,3,3,2,1,1,2,6,12,23,45,79,115,144,158,164,168,172,175,178,179,180,182,185,188,191,194,195,192,184,176,164,140,112,94,93,97,92,78,60,52,57,61,59,55,55,57,61,65,68,69,67,63,62,64,65,65,68,70,69,64,59,56,57,59,63,71,76,80,88,96,99,98,103,117,127,122,104,86,75,77,93,107,112,114,116,122,131,139,145,154,165,173,177,180,186,193,202,203,189,175,183,198,201,200,202,205,206,207,210,213,216,218,220,221,220,219,219,220,218,208,197,195,197,199,200,200,202,202,203,203,198,186,174,169,177,195,214,223,225,226,226,225,225,225,222,213,190,166,168,191,208,213,214,214,213,204,175,155,172,198,203,195,189,192,200,204,198,183,169,158,141,127,125,122,116,125,145,160,164,159,153,153,161,173,185,186,166,151,167,192,199,197,193,187,168,145,142,159,175,181,185,189,191,191,192,192,191,187,184,181,180,180,
29,24,13,4,2,3,9,24,50,80,99,96,80,73,83,96,111,133,156,170,175,176,175,174,165,136,86,40,17,9,5,3,2,2,3,3,4,4,4,4,5,5,5,4,3,2,1,1,1,2,4,9,23,46,75,110,141,157,160,161,162,166,169,172,175,179,183,185,186,188,189,186,180,172,159,141,123,115,121,130,128,110,86,73,80,86,79,72,76,87,100,107,109,104,92,78,68,66,67,69,71,74,76,76,72,69,66,66,72,84,97,107,119,134,144,149,154,162,165,155,139,125,113,114,134,155,163,165,169,174,180,185,186,187,189,191,194,197,203,208,211,208,193,183,194,211,217,217,218,220,220,219,219,221,223,225,226,226,225,222,219,217,216,213,211,212,215,215,213,211,211,213,216,217,216,211,207,206,210,217,222,222,221,222,223,222,220,220,220,210,180,144,139,165,191,204,209,207,202,193,169,152,167,187,188,176,170,177,189,195,192,184,178,177,172,166,161,151,143,157,178,189,191,189,187,187,190,195,198,190,165,147,164,189,197,196,194,186,158,119,105,129,160,177,184,187,187,187,188,190,190,188,186,185,183,182,
19,16,9,4,3,4,10,31,72,118,144,140,115,91,90,107,129,154,173,183,187,188,188,185,177,152,104,52,21,10,5,4,3,4,4,5,5,5,5,6,7,7,6,5,4,2,1,1,1,2,3,9,22,43,66,96,125,139,142,144,150,158,165,169,173,177,180,180,180,180,180,178,174,169,161,151,143,143,151,160,158,141,113,98,109,119,113,108,117,135,151,156,150,135,117,100,89,86,90,93,95,97,97,91,84,79,77,79,88,106,126,139,150,165,180,187,190,191,188,179,170,160,145,140,160,185,195,197,199,201,202,201,198,195,191,187,185,188,194,200,204,201,186,180,193,210,215,215,216,217,217,216,216,217,219,221,222,222,221,218,214,212,213,215,217,218,218,217,215,213,210,210,212,215,214,213,213,214,215,217,217,215,214,215,216,214,212,210,208,199,174,143,134,150,173,191,200,197,189,177,155,141,159,181,184,177,175,181,189,193,192,189,189,190,190,189,183,165,154,168,188,195,195,195,194,194,195,197,196,186,161,146,162,185,193,194,193,181,146,97,74,100,147,176,185,186,185,184,186,188,189,188,187,187,186,185,
9,8,5,4,8,14,24,50,95,142,168,168,147,124,121,135,152,169,182,187,189,188,186,181,170,148,105,54,21,10,7,6,6,6,7,7,6,6,7,8,9,9,8,7,5,4,3,3,5,7,10,14,27,46,68,95,121,133,136,140,149,161,168,172,176,180,182,182,182,182,182,181,180,180,179,176,173,174,180,184,182,166,137,120,136,156,157,155,161,173,182,184,173,157,143,135,130,129,133,137,139,139,133,119,105,97,97,102,114,134,154,168,177,186,196,201,201,197,188,179,172,163,145,138,160,186,197,199,202,204,203,200,195,189,183,177,174,175,178,184,193,191,175,167,182,197,199,202,207,209,209,210,210,210,211,212,213,213,212,210,207,205,208,211,213,214,213,211,210,209,206,205,206,208,208,208,207,207,208,207,207,206,206,206,207,206,204,203,202,197,185,171,162,162,169,183,192,192,186,172,145,131,153,182,190,188,189,192,194,194,192,192,192,192,192,192,185,165,151,165,186,193,192,192,192,192,193,193,191,183,163,151,165,184,191,192,189,170,128,79,60,91,144,178,187,185,183,182,184,187,188,188,188,188,187,187,
4,3,3,7,23,45,62,83,121,158,176,174,160,151,155,165,172,179,186,188,188,186,183,175,158,130,88,43,17,9,9,10,9,9,12,16,16,14,13,12,10,11,12,11,9,7,7,9,14,23,32,35,42,59,83,115,143,156,158,161,168,176,181,183,186,188,189,190,190,190,190,190,192,194,196,195,193,192,194,196,195,182,150,129,149,178,187,187,188,187,187,188,186,179,174,173,173,173,176,179,181,180,172,155,134,119,117,122,131,145,162,177,187,194,198,200,199,193,180,168,161,151,132,126,148,177,189,193,197,199,199,197,193,189,185,181,178,176,172,171,182,187,170,160,173,183,182,188,199,204,204,204,204,205,205,205,205,205,205,203,200,198,202,205,207,207,206,205,205,204,203,202,202,203,203,203,202,202,201,201,201,199,198,199,200,200,200,200,200,199,196,192,186,179,175,179,186,190,189,177,147,127,147,178,191,192,193,193,193,192,191,191,191,190,190,190,184,163,149,163,184,191,191,191,190,190,190,190,189,182,164,154,165,182,188,191,184,154,105,66,66,105,153,181,187,184,181,180,182,184,186,186,185,185,186,186,
2,2,3,14,44,83,104,116,142,168,178,169,157,158,170,179,182,182,181,177,174,174,171,160,138,103,61,28,12,9,12,15,14,17,28,42,46,38,26,19,16,16,16,15,14,14,15,18,29,50,70,72,67,79,107,143,170,182,185,186,188,190,192,193,194,195,196,196,197,197,196,196,198,200,201,200,197,196,197,199,198,186,152,128,149,183,197,198,195,185,178,185,195,198,197,197,197,198,199,201,202,201,195,180,154,131,128,135,140,147,161,177,189,195,197,199,198,194,185,176,171,161,139,128,150,179,190,193,196,197,196,196,195,194,193,191,189,185,173,165,176,185,173,162,171,176,171,178,193,201,201,201,200,201,201,201,201,201,201,199,193,190,194,200,201,201,201,201,200,200,200,200,199,199,199,199,199,199,199,200,199,195,191,193,197,198,198,198,198,197,197,196,194,188,181,177,180,185,189,181,151,127,140,169,185,189,190,191,191,189,189,190,190,189,188,189,184,167,155,167,184,191,192,192,191,190,190,189,188,181,161,149,158,174,182,185,174,140,95,74,91,132,167,185,188,185,182,180,181,182,182,178,176,176,178,179,
1,2,7,23,58,99,121,129,149,172,177,167,155,157,167,173,171,163,149,136,131,134,134,126,107,78,44,19,9,8,13,21,28,40,64,90,97,77,51,37,33,29,25,26,28,30,30,35,54,85,111,107,93,104,134,164,183,191,193,193,193,194,194,195,196,197,198,198,198,198,198,198,198,199,199,198,197,196,198,198,197,181,145,125,149,184,197,198,190,175,170,183,198,202,202,201,201,201,201,203,204,204,201,189,161,139,143,158,163,167,175,186,193,197,198,199,200,198,195,191,189,179,154,138,157,185,195,195,196,195,195,195,196,196,196,195,194,190,177,165,170,181,173,163,172,178,170,172,187,198,200,199,199,198,199,200,200,200,199,196,187,182,188,197,199,199,199,199,199,199,199,198,198,197,197,197,198,198,199,200,199,192,187,190,197,198,198,197,197,196,196,196,196,194,188,181,177,179,184,179,152,129,140,163,176,183,188,190,190,188,188,189,190,189,188,189,184,171,162,171,186,193,194,194,193,192,192,190,189,181,160,145,152,166,172,170,155,131,110,108,126,152,174,186,188,186,183,180,179,178,174,167,164,165,167,169,
1,2,9,26,54,84,105,120,143,167,173,164,153,147,143,138,131,117,97,79,79,93,103,100,91,78,54,27,11,9,17,31,50,77,110,139,145,122,88,69,60,49,43,47,57,64,66,73,93,122,139,127,113,129,159,177,185,189,191,191,191,191,192,193,195,196,196,197,197,197,197,197,197,196,196,196,195,196,197,197,192,171,134,121,151,185,196,194,181,167,168,184,197,200,199,198,197,197,197,198,199,200,199,191,167,150,161,180,186,189,192,195,197,198,198,198,199,199,197,196,195,186,159,142,160,187,196,196,195,194,194,195,196,196,196,196,196,194,184,168,167,175,168,158,171,183,174,168,181,196,200,199,199,198,199,200,201,201,200,196,184,176,184,196,199,199,199,200,200,199,199,199,198,198,198,198,198,199,199,200,198,190,185,190,197,199,198,198,198,198,199,199,199,198,195,189,181,177,179,175,151,133,146,166,171,174,183,188,190,189,189,190,190,190,189,189,184,169,160,171,186,193,194,195,195,194,193,191,189,182,164,146,148,157,156,144,132,130,136,144,148,156,169,182,186,184,181,177,175,172,167,161,160,160,159,159,
1,3,10,21,36,53,70,89,114,138,149,143,127,111,96,88,86,80,64,52,62,89,107,109,111,110,87,48,21,15,21,38,66,104,140,165,173,159,130,104,85,70,63,71,89,108,118,125,138,154,157,138,124,144,173,184,186,188,189,189,189,190,191,192,193,194,194,195,196,196,196,196,195,194,194,195,195,196,196,194,185,161,127,120,152,186,196,189,174,165,174,189,197,199,199,198,197,196,197,197,198,198,197,191,171,158,169,187,193,195,196,197,197,197,196,196,196,194,194,194,196,187,161,144,162,188,197,197,197,196,194,193,193,193,195,196,197,197,190,174,167,172,165,154,169,186,178,166,173,188,195,195,196,197,198,200,202,202,202,195,178,167,177,191,196,196,197,199,200,200,200,200,200,200,200,200,200,201,201,201,195,183,176,182,192,197,197,199,200,201,202,202,201,199,196,193,189,182,177,171,149,133,148,168,168,165,171,180,186,188,189,189,189,187,187,187,183,168,157,166,182,187,188,189,190,190,189,184,179,173,159,140,135,139,136,126,122,133,151,161,159,158,166,176,182,182,179,177,176,174,170,168,166,163,157,155,
3,6,15,26,31,32,38,51,71,92,102,97,81,64,56,61,72,76,70,63,74,99,118,128,141,143,113,64,32,25,28,38,64,105,143,168,179,176,158,131,106,90,85,91,110,136,157,168,174,178,172,146,128,149,178,188,189,189,188,186,184,184,186,189,191,193,194,195,196,197,197,196,195,195,196,197,197,198,197,191,176,153,129,125,154,185,192,180,165,166,181,194,198,199,200,200,199,199,200,200,200,199,199,191,169,154,166,186,194,196,197,197,197,197,196,195,191,186,184,189,195,189,162,144,162,191,201,200,200,197,192,186,182,184,189,193,195,198,194,180,172,176,168,156,171,190,184,167,163,171,177,181,186,190,193,197,201,202,202,193,169,152,161,176,180,179,183,188,193,195,198,199,200,201,201,200,200,200,200,200,191,171,157,163,178,186,190,193,196,198,199,200,199,195,192,191,191,188,181,171,149,132,142,159,160,153,154,163,174,181,184,184,182,179,177,181,183,170,156,159,168,169,166,167,170,171,166,156,147,141,133,121,119,127,132,134,137,146,160,169,171,170,170,174,180,184,184,184,184,183,182,181,178,171,163,160,
8,11,23,38,44,40,36,38,50,68,74,63,49,41,46,62,78,86,86,81,80,90,108,132,152,147,110,63,37,32,34,39,56,89,129,159,173,171,161,144,122,106,103,110,126,150,175,188,192,193,182,151,130,151,182,192,193,191,187,179,172,169,171,177,185,191,195,198,199,200,200,199,198,199,200,200,200,200,198,188,171,153,137,132,154,180,183,166,152,161,180,192,195,197,197,197,197,199,200,200,200,198,197,187,162,143,156,181,192,194,195,195,194,193,192,191,185,176,173,178,187,183,158,139,156,184,195,194,193,190,183,172,166,170,177,182,186,190,189,179,174,177,170,160,171,187,184,168,156,155,158,163,172,178,183,188,192,193,192,184,161,140,142,155,158,158,163,170,177,182,186,189,188,188,188,189,188,187,187,187,180,161,145,146,158,167,172,176,180,182,184,185,184,182,179,179,181,180,176,165,147,132,134,143,146,144,145,150,159,168,173,172,169,164,162,167,172,163,148,144,147,142,134,133,136,137,130,116,106,105,108,113,123,139,150,158,164,169,174,179,182,182,178,177,183,187,188,189,190,190,189,189,186,180,173,170,
16,17,23,36,48,57,60,58,65,84,87,67,48,44,51,62,73,79,84,84,76,71,87,116,134,124,89,54,36,33,34,35,46,72,110,144,155,148,143,139,123,106,108,124,142,160,175,185,189,190,179,149,130,149,177,188,188,185,178,168,158,152,153,161,173,183,189,192,195,196,196,196,196,196,197,196,195,194,190,179,167,158,148,141,153,170,171,156,146,154,169,177,180,182,181,180,182,184,186,188,187,184,180,173,152,137,147,167,177,180,180,179,176,173,174,175,170,162,157,159,164,160,142,128,140,161,169,168,165,162,157,151,146,148,152,155,159,163,163,159,159,162,158,153,158,166,166,156,147,144,144,147,153,159,162,165,167,167,166,161,148,132,127,135,141,141,144,148,153,157,161,162,159,156,157,160,160,158,157,159,156,147,137,135,138,143,146,148,150,151,152,153,154,153,153,153,153,153,152,146,136,128,128,131,134,139,143,143,144,149,153,151,147,143,141,143,145,139,129,128,129,122,114,114,118,120,116,106,102,110,123,136,151,165,174,180,184,187,187,188,189,189,186,184,187,189,188,189,191,191,191,190,189,185,182,180,
27,23,18,22,36,61,81,81,82,101,108,83,54,45,45,48,52,56,67,77,71,57,62,82,95,89,72,52,38,31,26,25,33,55,88,116,123,115,113,113,102,94,103,125,143,153,158,162,165,167,159,139,127,141,161,170,169,164,157,150,146,143,142,147,155,164,170,172,174,174,175,176,177,178,178,177,174,171,167,160,155,153,147,141,145,154,156,150,146,148,151,152,155,155,153,153,156,159,161,163,162,158,154,152,144,137,141,150,155,155,155,153,148,145,148,150,148,143,140,138,137,134,126,119,124,135,139,138,134,131,130,129,127,127,126,126,130,133,134,135,138,141,141,139,139,141,142,139,136,135,135,135,138,140,141,142,142,142,142,141,137,128,123,127,132,133,133,133,135,136,138,137,133,128,130,134,135,135,135,135,135,131,127,124,122,122,122,122,123,124,124,125,126,128,130,131,131,132,133,132,128,126,126,127,129,135,140,137,134,137,140,139,136,134,133,130,127,124,123,129,133,127,124,130,137,142,143,140,141,151,163,172,179,185,189,191,193,193,192,191,192,193,191,189,190,191,190,190,190,190,189,189,189,188,188,188,
38,31,18,14,28,60,88,89,81,94,104,84,53,37,34,33,32,35,48,64,64,50,44,52,58,62,63,55,42,31,21,17,21,40,65,81,84,81,79,77,76,85,104,123,135,139,140,142,144,146,144,136,131,137,148,153,152,146,138,136,140,142,141,141,145,150,153,154,154,154,154,155,156,156,157,155,152,148,146,143,142,141,136,133,135,140,143,142,143,143,141,139,142,144,144,145,148,151,152,153,153,150,148,149,149,148,149,151,151,150,149,148,145,143,145,148,147,146,145,143,141,140,138,135,136,139,141,141,139,137,136,137,137,136,134,133,136,139,140,141,145,148,149,148,147,148,148,147,146,146,147,147,148,148,149,149,150,150,150,150,149,146,144,145,147,147,147,146,146,146,147,146,142,139,140,144,145,146,146,145,143,140,137,133,130,128,127,128,128,129,129,130,132,136,140,142,143,144,146,146,145,143,143,144,144,147,149,148,148,151,156,157,157,157,156,153,149,147,149,155,160,158,158,164,171,175,178,178,179,184,188,190,191,193,194,194,194,194,192,191,192,194,193,192,193,193,193,192,191,188,187,187,189,190,191,191,
51,41,21,15,34,71,97,92,74,74,83,75,52,39,39,39,34,32,40,52,54,47,41,41,42,44,49,47,38,29,22,18,20,33,50,60,62,62,59,55,66,91,118,134,142,147,150,151,152,154,155,154,152,152,156,159,159,154,148,148,153,157,157,157,158,160,159,156,156,158,159,159,159,159,159,158,155,152,150,150,151,148,143,142,145,149,150,151,153,155,155,156,160,164,166,168,171,173,173,174,174,173,172,173,174,174,174,175,174,174,174,174,173,172,174,175,175,176,176,175,174,173,173,172,171,172,173,173,173,172,172,172,172,172,171,170,172,173,174,176,177,179,179,179,179,180,180,179,178,178,178,179,179,179,180,180,181,182,182,181,180,179,179,179,180,180,180,179,179,179,179,179,177,175,176,178,178,179,178,177,175,172,169,166,163,161,160,161,161,161,162,162,165,170,174,175,176,176,177,177,176,175,175,176,175,175,175,176,178,181,184,186,187,187,187,185,183,182,182,184,186,185,185,188,190,192,192,192,193,194,194,194,193,194,195,195,195,194,193,191,192,193,194,194,194,194,195,194,193,190,187,187,189,191,191,191,
60,47,24,17,41,81,104,92,65,53,60,61,51,47,56,62,57,50,48,50,48,44,42,40,35,30,30,30,27,25,26,28,31,37,45,52,56,54,49,48,67,104,134,149,160,169,175,177,178,178,179,180,179,178,178,179,180,178,176,175,178,181,181,181,181,180,177,172,173,177,179,179,179,180,179,178,175,169,165,168,173,171,166,167,172,174,174,176,179,182,182,184,187,190,192,194,196,197,197,197,197,198,198,197,196,196,197,197,197,197,198,198,198,198,198,199,199,199,199,199,198,198,198,198,197,197,197,197,197,197,197,197,197,197,197,197,197,198,199,199,200,200,200,200,201,201,201,200,200,200,200,200,201,201,201,201,202,202,202,201,200,200,200,200,201,201,201,201,200,200,200,200,200,199,200,200,200,200,199,198,197,195,194,192,190,189,189,189,188,188,189,190,192,194,196,197,197,197,196,196,196,195,195,195,195,195,195,195,196,197,198,198,199,199,198,198,197,196,196,195,195,195,195,195,196,196,196,196,196,196,195,195,194,195,196,196,195,195,195,194,194,195,195,196,196,196,196,196,195,193,191,190,191,191,191,191,
53,43,24,17,35,67,83,71,47,34,37,43,43,48,65,78,78,72,66,62,54,43,37,33,27,21,19,20,21,24,32,41,46,45,44,44,43,39,34,37,63,101,129,145,162,179,188,191,191,191,191,192,192,192,192,192,193,192,192,192,193,194,194,194,193,192,188,185,186,189,190,191,191,192,192,190,184,174,168,174,183,181,178,180,185,187,189,194,197,198,198,199,200,201,201,202,203,203,203,204,204,204,204,203,202,202,203,203,203,204,204,204,203,203,204,204,204,204,204,204,203,203,203,203,203,203,202,202,202,202,202,202,202,202,202,202,202,203,203,204,204,204,204,204,205,205,204,204,204,204,204,204,204,204,204,205,206,206,206,205,204,204,203,203,204,205,205,205,204,204,204,204,204,204,204,204,204,203,203,203,202,202,201,201,200,199,199,199,198,198,198,199,200,201,200,200,200,201,201,201,200,200,200,199,199,200,200,200,200,199,199,200,200,200,199,199,199,198,198,198,197,197,197,197,198,198,198,198,197,197,197,197,197,197,197,197,197,197,197,197,197,197,197,198,198,198,198,197,197,196,195,194,194,193,193,193,
33,29,19,13,20,35,42,36,26,19,20,24,30,43,61,75,80,79,76,73,61,44,30,22,17,16,18,21,24,31,44,58,61,54,46,38,30,27,24,30,55,87,108,125,152,177,190,192,192,192,193,193,194,195,195,195,195,195,195,195,195,196,196,196,195,195,194,192,192,192,192,192,192,193,192,187,178,168,166,173,180,180,178,179,180,183,191,198,201,202,202,202,202,202,202,202,202,202,203,203,203,204,204,203,202,202,203,203,203,203,203,202,201,202,203,203,203,203,203,203,203,203,203,202,202,202,202,201,201,202,202,202,202,203,202,202,202,202,203,204,204,204,204,204,204,205,204,204,204,204,205,204,204,203,203,204,204,205,205,205,204,203,203,202,203,204,204,204,203,203,203,203,203,203,203,203,203,203,202,202,202,202,202,202,202,201,201,201,200,200,200,201,201,200,200,199,200,201,202,201,201,201,200,200,200,200,201,201,200,200,200,200,201,201,200,200,200,199,199,199,199,199,199,199,200,200,200,200,199,199,199,199,200,199,199,199,199,199,199,199,198,199,199,199,199,199,199,199,199,198,198,198,197,196,196,195,
14,15,13,11,11,14,14,12,11,10,10,13,21,35,51,61,69,76,77,70,57,42,27,16,12,13,19,26,32,45,66,82,81,71,59,44,34,37,40,43,60,85,101,120,151,179,191,193,192,192,193,193,194,195,195,195,195,196,195,195,195,195,196,196,196,196,197,196,195,194,193,192,192,192,190,184,173,166,168,173,176,177,179,179,178,181,191,199,201,202,202,202,202,202,202,202,202,202,202,202,203,203,204,203,202,202,203,203,203,203,202,201,201,201,203,203,203,202,202,202,202,201,201,201,202,202,201,201,201,202,202,202,202,203,203,202,202,202,203,204,204,204,204,204,204,205,204,204,204,204,204,204,204,203,203,203,203,204,205,205,204,203,203,202,202,203,203,203,202,202,202,202,202,202,202,202,202,203,203,202,202,202,202,202,202,202,202,201,201,201,201,201,201,200,200,200,201,202,202,201,201,201,201,201,201,201,201,201,201,200,200,201,201,201,200,200,200,200,200,200,200,199,199,199,199,200,200,200,199,199,199,200,201,201,200,200,200,200,199,199,198,199,199,199,199,198,198,198,198,198,198,198,198,198,197,196,
6,8,10,9,9,8,6,5,6,7,8,9,15,28,42,48,60,78,81,66,49,37,26,15,10,12,17,26,40,61,90,110,111,99,82,61,51,63,78,81,89,107,121,137,163,184,192,193,193,193,193,194,194,195,195,195,195,195,195,194,194,194,195,195,196,196,197,197,196,195,194,193,193,193,192,187,178,174,176,178,178,180,184,185,185,188,195,199,200,200,200,200,200,200,200,200,200,201,201,201,201,202,202,202,201,201,202,202,202,202,201,201,200,201,202,202,202,201,201,201,200,200,200,200,201,201,201,200,200,200,200,201,201,201,202,202,202,202,202,203,203,203,203,203,203,203,203,203,202,202,202,203,203,202,202,202,202,203,203,204,203,202,202,201,201,201,201,201,201,200,200,201,201,200,199,200,201,201,202,201,201,200,201,201,201,201,201,201,201,201,201,201,200,200,200,200,201,201,200,200,200,200,200,200,200,200,200,200,200,199,199,200,200,199,199,199,199,199,199,198,198,197,196,196,196,197,197,197,197,197,197,198,199,198,197,197,197,196,196,196,196,196,197,197,196,196,195,195,195,196,196,196,196,196,195,195,
4,5,6,7,6,5,4,4,5,5,6,8,13,24,35,43,59,82,88,69,46,32,21,14,10,11,14,23,45,75,109,134,140,127,104,79,68,85,113,126,129,135,144,157,175,187,191,192,192,192,192,192,193,193,193,193,193,193,193,193,193,193,193,194,194,194,195,195,194,194,193,193,193,193,193,191,188,186,187,186,186,188,190,192,193,195,197,198,198,198,197,197,197,197,197,197,198,198,198,198,198,199,199,199,199,199,199,200,200,199,199,199,199,199,199,199,199,199,199,199,198,198,198,198,199,199,199,198,198,198,198,198,198,198,198,199,199,200,200,200,200,200,200,200,200,200,200,200,199,199,199,200,200,200,199,199,200,200,200,200,200,199,198,198,198,198,197,197,197,198,198,198,198,197,197,197,198,198,199,198,198,198,198,198,198,198,198,198,198,198,198,198,198,198,198,197,197,197,196,196,197,197,197,196,196,196,196,196,196,196,196,196,196,195,195,194,195,195,195,194,194,193,192,192,191,192,192,193,193,193,192,193,193,193,192,192,191,191,191,191,191,191,191,191,191,191,191,190,191,191,191,191,191,191,191,191,
3,3,3,4,3,3,3,4,5,5,5,8,14,21,28,38,57,77,81,67,45,27,16,11,11,11,14,24,49,86,123,152,161,145,114,88,80,96,127,152,159,158,160,170,181,187,188,189,189,189,189,189,189,190,190,190,190,190,190,190,190,190,190,191,191,191,191,191,191,190,191,191,191,190,191,191,191,191,191,191,191,192,193,193,194,195,195,195,194,194,194,194,194,193,193,194,194,194,195,195,195,195,195,195,195,196,196,196,195,195,195,195,195,195,195,195,195,195,195,195,195,195,194,195,195,196,196,195,194,194,194,194,194,194,194,194,195,196,196,196,195,195,194,195,195,196,196,195,195,195,196,196,196,195,195,195,195,195,195,195,194,193,193,193,193,193,193,193,193,194,194,195,194,194,193,194,194,194,195,195,195,194,194,194,194,194,194,193,193,193,193,194,194,193,193,192,192,192,192,192,193,193,192,191,190,190,190,191,192,192,191,191,190,190,189,189,189,190,190,189,189,190,190,189,189,189,189,190,190,190,189,189,188,188,187,186,186,185,185,185,185,185,185,185,186,186,186,186,186,186,187,187,186,187,187,187,
3,2,2,2,2,3,3,4,5,5,6,10,18,22,23,30,46,56,56,48,35,21,12,10,13,16,20,28,52,89,129,159,168,150,116,92,88,101,127,156,173,174,174,177,182,184,184,185,185,185,185,185,185,185,185,186,186,187,187,187,187,187,187,188,188,188,189,188,188,187,187,187,187,187,187,187,187,188,188,188,189,191,191,192,192,193,192,192,191,191,190,190,190,189,189,190,190,190,191,191,191,191,192,193,193,193,193,193,192,192,193,192,192,191,191,191,191,191,191,191,190,190,191,192,193,193,193,193,192,192,192,192,192,192,192,192,192,192,192,192,191,190,189,190,191,191,191,191,191,192,192,192,192,191,191,191,191,191,191,190,189,189,189,189,188,189,189,189,189,189,190,190,191,191,190,190,191,192,192,192,192,191,191,191,190,189,188,188,188,188,188,188,188,187,187,187,188,189,190,190,190,190,188,186,185,186,186,188,189,189,187,186,185,185,184,184,184,185,185,185,186,188,189,190,189,189,190,190,190,190,189,189,189,188,185,183,181,181,180,180,180,180,180,181,182,183,185,185,185,185,186,186,186,186,186,186,
3,3,3,2,2,3,4,4,5,6,8,13,22,26,22,21,27,31,28,24,20,13,8,9,15,21,26,33,52,85,123,154,165,152,122,103,103,112,130,156,175,180,180,180,181,181,181,181,181,181,181,181,181,181,181,182,184,185,186,186,186,187,187,188,188,189,189,189,188,186,184,184,183,184,184,184,184,184,184,185,187,190,192,192,192,193,193,192,191,190,188,187,186,186,186,187,188,187,187,187,187,189,192,193,194,194,194,193,193,193,194,193,192,189,188,188,188,188,188,187,186,186,187,189,192,194,195,195,195,194,194,194,194,194,194,193,192,191,190,189,188,187,186,187,188,188,188,188,189,189,189,189,189,188,188,188,187,187,188,187,187,186,186,186,186,186,186,187,186,186,186,186,187,188,188,187,188,188,189,189,189,189,189,189,187,185,183,183,183,183,183,183,183,182,182,182,184,186,187,187,187,186,184,183,182,183,183,184,185,185,183,181,180,180,180,180,180,181,181,181,183,186,188,188,188,188,188,188,188,188,188,188,188,187,184,180,178,177,177,177,177,177,178,178,179,181,183,185,184,184,184,184,185,185,185,185,
3,3,4,3,2,3,3,3,4,6,10,15,23,26,20,14,14,15,13,10,9,7,6,7,13,20,26,34,50,77,112,142,158,152,134,124,127,133,143,161,175,179,179,179,178,178,178,178,179,179,178,178,177,177,178,179,181,184,186,186,186,187,187,188,189,189,190,189,187,184,182,180,180,180,181,181,181,181,181,182,184,188,191,192,192,192,192,191,191,189,186,184,183,183,183,184,185,185,184,184,185,187,190,193,194,195,194,194,193,194,194,194,191,188,186,185,186,186,186,185,184,184,185,187,191,194,197,197,197,196,195,194,194,194,194,193,191,189,187,186,185,184,184,185,185,186,186,185,186,187,187,187,186,186,186,186,185,185,186,186,185,184,184,184,184,184,185,185,184,184,183,183,184,184,184,184,184,184,185,185,185,185,185,184,183,181,180,180,180,180,179,179,179,179,179,180,180,181,181,181,180,179,178,178,178,178,178,178,178,178,177,175,175,176,176,176,176,177,177,178,179,180,182,182,181,181,181,181,181,181,181,182,182,181,179,176,174,174,174,174,174,174,174,175,175,177,178,179,178,177,177,177,177,178,178,178,
3,3,3,3,2,2,2,2,3,6,10,17,21,21,14,8,8,9,7,5,5,4,4,6,10,15,21,31,46,73,106,135,151,150,141,140,148,154,159,168,175,176,176,176,175,175,176,176,177,177,176,175,174,174,175,176,178,180,181,182,182,182,182,183,184,185,185,184,183,180,178,177,177,177,177,178,179,179,179,179,180,183,185,186,186,186,185,185,186,185,183,182,181,180,181,182,182,182,182,182,182,184,186,187,188,189,189,188,188,189,189,189,187,184,183,183,183,183,183,183,182,182,183,184,187,189,191,192,191,190,188,188,188,188,189,188,187,184,183,183,182,182,182,182,182,182,182,182,183,184,184,184,184,184,184,183,183,183,184,184,183,182,182,182,182,182,182,182,182,182,182,181,181,181,181,181,181,180,181,181,182,182,181,180,179,179,178,177,178,177,176,176,176,177,177,177,177,177,176,176,175,175,174,174,174,174,174,173,173,173,172,172,172,172,172,172,172,173,173,174,174,174,175,174,173,173,173,173,173,173,173,174,174,173,172,171,170,170,170,170,170,169,169,169,170,170,171,171,170,169,169,168,168,168,169,169,
2,2,2,2,2,2,2,2,3,4,9,14,17,14,8,5,5,5,5,3,3,3,3,5,8,12,16,25,42,70,103,131,146,147,144,149,158,163,167,171,174,174,173,173,173,173,173,174,174,174,173,173,172,171,172,173,174,174,175,175,175,175,175,175,176,178,178,178,177,176,175,174,174,174,175,175,176,177,177,177,177,177,178,179,179,179,179,179,180,180,180,179,178,178,178,179,180,180,180,179,179,180,181,181,181,181,181,181,181,182,182,183,182,181,180,180,181,181,181,180,179,180,181,181,182,183,184,184,184,182,180,180,180,181,182,182,181,180,180,180,180,179,179,179,179,179,179,179,180,181,181,181,181,182,181,180,180,180,181,181,180,180,180,180,179,179,179,179,179,179,179,179,179,179,179,179,178,178,178,178,179,179,178,177,177,176,175,175,175,175,174,174,174,175,175,175,175,175,174,173,173,172,172,172,172,172,172,171,171,171,170,170,169,169,169,169,169,170,170,170,169,169,170,169,168,168,168,168,168,168,168,168,168,167,166,166,166,166,166,166,165,164,165,164,164,164,165,165,164,164,164,163,162,162,162,163,
1,1,1,1,1,1,2,2,2,3,6,10,12,10,6,3,3,3,2,2,2,2,2,4,6,8,11,20,38,65,97,124,139,144,150,158,164,166,168,170,171,171,171,170,170,170,170,170,171,171,171,170,169,169,169,170,171,171,171,171,171,171,171,171,172,174,174,174,173,172,172,172,173,173,173,173,174,175,175,174,174,174,174,175,175,175,175,175,176,177,176,176,176,175,175,176,177,177,177,177,177,177,177,177,177,176,177,177,177,178,179,179,179,179,179,178,178,178,178,178,177,177,177,178,179,178,178,178,178,177,176,175,176,177,177,177,178,178,178,178,178,177,177,177,177,176,177,178,179,180,179,179,179,180,179,178,178,178,179,179,179,179,179,178,177,177,176,176,176,177,177,177,176,176,176,176,176,176,175,176,177,177,176,175,175,174,174,173,173,173,173,172,173,173,173,173,173,173,173,172,171,171,170,171,171,171,170,169,169,169,168,168,167,167,167,167,168,168,168,167,166,166,166,166,166,166,165,165,165,165,165,165,165,164,164,164,164,164,164,163,162,162,161,161,160,160,161,161,161,161,161,161,159,159,159,159,
1,1,1,1,1,1,1,1,1,2,4,7,9,8,5,3,2,2,1,1,1,1,1,3,4,5,8,17,34,60,90,117,133,144,156,166,168,167,167,168,169,169,169,168,168,168,168,168,168,168,168,167,167,167,168,169,170,170,169,169,169,169,170,170,171,172,172,171,170,170,170,170,171,172,172,171,172,172,172,171,171,171,171,172,173,173,173,172,173,173,173,173,173,172,172,173,174,175,174,174,174,174,174,174,174,174,175,175,175,176,176,177,177,177,177,176,175,175,176,176,175,174,174,175,176,175,174,174,174,174,173,172,173,174,174,174,175,175,175,176,175,175,174,175,175,175,175,176,177,177,177,176,177,178,178,177,177,177,176,176,177,177,176,176,175,175,174,174,174,175,175,174,174,174,174,174,174,174,174,174,174,174,173,173,173,172,172,172,172,172,171,171,171,171,171,171,171,171,171,171,170,170,170,170,170,169,168,168,168,168,168,167,167,167,167,167,167,168,167,165,164,164,165,165,165,165,164,164,164,164,164,164,163,163,163,163,163,163,163,162,161,160,160,159,158,157,158,158,158,159,160,160,158,158,157,157,
1,1,1,1,1,1,1,1,2,2,4,6,7,6,4,2,2,1,1,1,1,1,1,2,3,4,7,16,35,62,90,112,128,146,161,169,169,168,168,168,168,168,168,167,166,166,166,167,167,166,165,165,166,167,167,168,169,169,169,168,168,169,170,171,171,171,170,169,169,169,169,169,169,170,170,170,170,169,169,169,169,169,169,170,171,171,171,170,170,170,170,171,170,170,170,170,172,172,172,172,171,171,171,172,172,172,173,173,173,173,174,175,175,174,174,173,172,172,173,173,173,172,172,173,173,172,171,170,171,171,171,171,172,172,172,172,173,173,173,173,173,172,172,173,173,173,174,174,174,174,174,174,175,175,176,175,175,174,174,174,174,174,174,174,173,172,171,171,172,173,173,172,172,173,173,173,173,173,173,173,172,171,171,172,172,172,172,172,172,172,172,171,171,171,170,170,170,171,171,170,170,171,171,171,170,169,167,168,169,169,169,169,168,168,168,168,169,169,168,166,165,166,166,166,165,165,165,165,165,165,165,164,163,163,163,164,164,164,164,164,163,162,161,160,158,157,157,158,159,160,160,160,159,159,159,159,
1,1,1,1,1,1,2,2,2,3,4,5,5,4,2,1,1,1,0,0,1,1,1,2,3,4,10,25,51,81,100,110,127,150,165,170,169,169,169,168,168,168,167,166,165,165,166,166,166,165,165,165,166,166,167,168,169,169,169,168,168,169,170,171,170,170,169,168,168,169,169,168,168,168,169,170,169,168,168,168,168,168,169,170,171,171,170,169,169,169,169,170,170,169,169,169,171,172,172,171,170,169,169,170,171,171,172,172,172,172,173,173,173,172,172,172,172,172,172,172,172,172,172,172,172,171,170,169,170,171,171,171,172,172,172,172,172,172,171,171,172,172,172,172,172,172,172,172,172,172,173,173,173,173,173,174,173,173,173,173,173,173,174,174,172,171,170,170,171,173,173,173,174,174,174,174,174,174,174,173,173,173,172,173,173,173,173,174,174,175,174,173,173,172,172,173,172,172,172,172,172,173,173,172,171,169,168,169,171,172,172,171,171,171,170,171,171,171,171,170,169,169,169,169,167,167,168,168,168,168,167,166,166,165,166,166,166,167,168,168,167,166,165,164,162,160,160,161,163,163,163,162,162,162,162,162,
2,2,1,1,1,1,2,2,2,3,3,3,3,2,1,1,1,0,0,0,1,1,1,2,4,9,21,45,77,102,111,118,136,157,168,169,169,169,170,169,169,168,168,167,166,166,167,166,166,166,167,167,167,167,168,168,169,169,169,169,169,170,170,171,170,169,169,169,169,170,170,170,168,168,169,170,170,170,170,170,170,170,171,171,171,172,171,170,169,170,171,171,171,170,170,171,172,173,173,171,170,169,169,170,172,172,173,173,173,173,173,173,173,173,173,173,174,174,174,174,174,175,174,174,174,173,172,172,172,173,173,173,172,172,173,174,174,174,173,173,173,173,173,174,174,173,173,173,173,174,175,175,174,174,174,174,174,174,174,174,174,175,176,176,174,173,172,172,174,175,175,176,176,176,176,176,175,176,175,176,176,177,176,175,175,175,175,176,177,177,177,176,175,175,175,175,175,174,173,173,174,175,175,173,171,170,170,171,173,174,174,174,174,174,173,173,173,174,174,174,173,172,172,172,171,171,171,171,171,171,170,169,169,168,169,169,170,171,171,171,171,170,169,168,166,165,165,167,167,167,166,165,165,165,165,165,
3,3,2,1,1,1,2,2,2,2,2,1,1,1,1,0,0,0,0,0,1,1,2,4,9,20,39,65,92,112,123,136,154,166,169,169,169,170,170,169,169,169,168,168,168,168,168,168,168,168,169,169,169,169,169,169,169,170,170,170,170,171,171,171,171,170,170,170,171,172,172,172,171,170,171,172,172,172,173,174,174,173,173,173,173,173,173,172,172,173,173,173,173,172,173,174,175,175,174,173,173,172,172,174,175,175,176,176,175,175,175,175,175,175,175,176,177,177,177,177,177,178,178,177,177,176,176,175,176,176,175,175,174,174,175,176,177,177,176,175,175,176,176,176,176,176,176,175,176,177,178,179,178,178,177,177,177,176,177,177,177,177,178,178,177,176,175,176,177,178,178,177,177,177,177,177,176,176,176,177,179,180,179,178,177,177,176,176,177,178,178,177,177,177,177,177,176,175,174,174,174,175,175,174,173,172,172,173,174,175,175,176,176,175,174,174,174,175,176,177,176,175,174,174,173,173,173,173,173,172,172,172,171,170,170,171,172,172,172,172,172,172,171,170,169,169,169,170,170,168,167,166,167,167,167,166,
5,4,2,1,1,1,1,2,1,1,1,1,1,1,0,0,0,0,0,1,1,3,5,8,16,32,54,77,101,122,140,156,167,170,170,170,169,169,169,169,169,169,169,169,170,170,169,169,169,169,169,169,169,169,169,169,169,170,171,171,172,171,171,171,171,170,170,171,172,172,173,173,173,173,173,173,173,173,174,176,176,175,174,174,174,174,173,173,173,175,175,175,174,174,175,176,176,175,175,174,175,175,176,177,178,177,177,176,177,177,177,177,176,176,176,177,178,178,177,178,178,179,179,179,179,178,178,178,178,178,177,176,176,176,177,177,178,178,178,177,177,178,178,178,178,178,178,177,178,179,180,181,182,181,181,180,179,179,179,179,179,179,179,179,178,177,177,177,178,179,179,178,177,176,177,176,176,176,176,177,178,180,179,178,178,177,177,176,177,177,177,177,178,178,177,177,176,175,174,174,174,175,175,175,174,173,173,174,175,176,176,176,176,175,173,174,174,175,177,178,178,176,174,174,174,174,174,174,174,173,173,173,172,171,170,171,172,172,171,171,171,171,171,170,170,170,170,171,170,169,168,168,168,168,167,167,
7,6,3,2,1,2,2,2,1,0,0,0,0,0,0,0,0,0,1,1,2,5,10,14,22,39,62,88,114,136,153,165,170,171,170,169,169,168,168,168,169,169,169,170,171,170,169,169,169,169,168,169,169,168,168,168,169,169,170,171,172,171,171,170,170,170,170,171,172,172,172,173,173,174,173,173,172,172,174,175,176,175,175,174,174,174,174,174,174,175,176,176,175,175,175,176,175,174,174,174,175,177,178,178,178,177,176,175,176,177,177,177,177,177,178,178,178,178,177,177,178,179,179,179,179,179,179,179,179,178,177,177,178,178,179,179,179,179,179,178,178,179,179,178,178,179,178,178,179,180,180,181,182,182,182,181,181,180,180,180,180,180,180,180,179,178,177,178,179,180,179,178,177,177,177,177,176,176,176,176,177,178,178,177,177,178,177,177,176,176,177,178,178,178,177,176,176,176,175,175,175,175,175,175,175,175,175,175,175,176,176,176,176,175,174,175,175,175,176,177,177,175,174,175,175,175,175,175,175,174,174,173,173,173,172,172,172,172,171,171,171,171,171,170,170,169,170,171,171,171,170,169,169,168,167,167,
10,8,4,2,2,3,4,2,1,1,1,1,1,1,0,0,0,0,1,1,3,8,15,21,28,44,72,102,125,142,155,165,170,171,170,169,169,168,168,168,169,170,170,171,171,170,169,169,169,169,169,168,167,166,166,168,169,170,170,171,171,171,171,171,171,171,171,171,171,171,172,172,173,174,174,173,173,172,174,175,176,176,176,175,174,175,176,176,175,175,176,176,176,176,176,176,175,174,174,175,176,178,179,179,178,177,176,176,176,177,178,178,179,179,179,179,179,178,178,178,179,179,179,179,180,179,179,179,180,179,178,178,179,180,180,180,180,180,179,179,179,179,179,179,179,179,179,179,179,179,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,179,179,179,180,181,181,180,179,179,179,178,177,176,177,178,179,178,178,177,177,177,177,177,177,177,178,178,179,178,178,177,177,177,177,176,176,175,175,176,176,176,176,176,176,177,177,177,177,176,176,176,176,176,176,176,176,175,175,175,176,176,176,177,177,176,175,174,174,174,174,173,173,173,173,173,173,172,172,172,171,171,172,172,173,173,172,171,170,169,169,169,
11,9,5,3,3,4,4,3,2,2,2,2,2,2,1,1,1,1,1,1,3,10,25,40,48,60,87,114,130,140,152,164,171,172,172,171,171,171,170,170,170,171,172,172,172,171,170,170,170,169,168,166,162,159,162,168,171,172,172,173,173,173,172,172,173,174,174,173,173,173,174,174,175,176,176,175,175,175,176,177,178,178,178,177,175,176,177,178,178,178,178,178,178,177,177,177,177,177,177,178,179,180,180,180,179,179,178,178,178,179,180,180,180,180,180,181,180,179,179,180,180,180,179,180,180,180,180,180,181,181,180,180,180,181,181,181,181,181,181,181,181,181,181,181,181,181,181,180,180,180,180,180,181,181,180,179,180,181,182,182,182,182,183,184,183,181,180,181,181,182,183,182,182,181,181,180,179,177,179,181,181,180,179,178,178,176,176,177,179,180,180,180,179,179,179,179,178,178,178,178,177,177,177,177,178,178,179,179,180,180,180,180,180,180,180,179,179,178,178,178,178,177,177,178,179,179,179,179,179,179,178,177,177,177,177,177,177,177,176,176,176,176,176,176,176,176,176,176,175,175,174,173,172,172,172,172,
9,7,4,3,3,4,3,3,3,5,6,7,6,4,3,3,3,2,2,3,6,19,44,71,80,83,99,122,136,144,155,167,173,174,174,174,174,174,174,173,173,174,175,175,174,172,171,171,169,165,159,154,147,143,149,163,173,175,176,177,177,177,176,176,177,178,178,178,178,179,179,179,179,179,178,178,178,178,179,180,180,180,180,180,178,177,178,179,180,180,180,181,180,180,180,180,180,180,181,181,181,182,182,182,181,181,181,181,181,181,182,182,182,182,182,183,183,182,183,183,184,183,182,182,183,183,182,183,183,183,183,182,181,182,183,183,183,183,182,182,183,183,184,184,184,184,184,184,183,183,182,182,183,183,181,180,181,183,184,184,183,183,184,185,185,183,183,183,183,184,185,184,183,183,183,182,181,180,181,183,183,182,180,180,180,178,177,179,181,182,182,182,181,180,180,180,180,180,180,180,180,179,179,180,181,183,184,185,186,185,185,185,185,185,185,185,184,184,184,184,183,182,182,183,184,185,185,184,184,183,183,182,182,183,184,183,182,182,181,181,181,181,181,181,182,182,181,180,178,177,177,176,175,174,174,174,
6,5,3,3,3,4,5,5,6,8,11,12,10,6,4,5,5,5,7,10,15,29,57,85,93,93,105,127,145,156,165,172,176,177,176,176,177,177,177,177,177,178,179,179,177,175,174,173,167,152,137,128,122,120,131,155,174,181,182,183,183,183,183,183,184,184,184,184,185,186,186,186,185,183,181,180,180,181,181,182,182,181,181,181,180,179,180,181,181,182,182,183,183,183,182,182,183,183,184,183,183,184,184,184,184,183,183,182,183,183,184,184,184,184,184,185,186,187,189,189,190,189,188,188,189,189,188,188,189,188,187,185,185,185,185,186,186,185,185,186,186,187,187,187,187,187,188,187,187,187,186,186,187,186,185,183,184,186,186,186,185,185,186,186,185,184,184,185,185,186,186,185,185,185,185,185,184,184,185,185,184,183,183,183,184,183,181,182,184,184,183,183,182,181,181,182,182,182,182,182,182,181,182,182,184,186,188,189,189,188,188,188,189,189,188,188,187,188,189,189,188,186,185,186,187,187,187,187,187,186,186,186,186,187,187,187,186,185,185,184,184,184,184,184,184,184,184,182,180,179,178,177,176,175,175,174,
4,4,3,2,3,5,8,10,10,10,12,13,10,7,7,9,10,12,16,21,24,34,54,72,81,90,107,130,151,165,173,176,178,178,178,177,178,179,180,181,181,182,182,183,182,181,180,177,163,135,107,97,99,104,117,145,172,183,186,186,187,187,187,187,187,188,188,188,188,189,189,189,188,186,183,181,181,182,182,182,182,181,181,181,181,181,181,181,182,182,183,183,184,183,183,184,185,185,185,184,184,184,185,185,185,185,184,184,184,185,186,185,185,185,185,186,187,190,192,193,194,194,193,193,194,193,192,192,192,192,190,188,187,187,187,188,188,187,188,188,189,189,188,188,188,189,189,189,189,189,189,189,189,189,188,186,186,187,188,188,187,187,186,186,185,184,184,186,187,187,187,186,186,187,187,187,187,187,187,185,184,185,186,186,186,186,185,185,185,184,184,183,182,182,182,182,182,182,182,183,183,183,183,183,184,184,185,185,185,185,185,185,185,186,185,185,185,185,186,187,186,184,182,183,183,183,183,183,183,183,183,183,183,183,183,183,183,183,182,182,182,181,181,180,180,181,180,179,178,177,177,176,175,174,173,173,
4,4,3,2,2,5,11,15,14,11,10,10,10,11,14,18,22,28,34,35,33,36,45,54,66,86,111,134,154,168,176,177,178,178,178,178,177,178,179,181,182,182,183,183,184,183,182,178,159,120,83,73,85,95,108,135,165,180,183,184,184,184,184,184,184,184,184,184,185,185,185,185,185,183,181,181,181,181,181,181,181,180,180,180,180,181,181,181,181,181,182,183,183,182,182,184,185,184,184,184,184,183,184,185,185,185,184,184,184,185,185,185,184,185,185,185,186,188,190,191,191,191,191,191,192,191,190,189,190,190,189,187,186,186,186,186,186,186,186,188,188,187,186,186,186,186,187,187,187,188,188,189,189,188,187,187,187,187,187,187,187,186,186,186,185,184,184,185,186,187,186,186,187,187,188,187,186,187,187,186,185,185,186,186,186,185,185,184,184,183,183,182,181,181,182,181,180,181,182,182,182,182,182,182,181,181,181,180,179,179,180,180,180,181,181,180,180,180,181,181,180,178,177,177,177,177,177,177,178,178,178,177,177,177,177,178,177,177,177,177,176,176,175,174,173,174,173,173,172,173,172,172,172,171,171,171,
4,4,3,2,2,5,12,17,17,13,10,10,14,21,27,30,37,47,55,54,45,39,37,42,55,82,114,141,160,171,176,176,176,178,178,178,177,176,176,178,179,179,179,180,181,181,180,173,151,108,67,57,70,82,100,131,161,175,178,179,180,179,179,178,178,179,179,179,179,179,180,180,180,179,179,180,180,180,180,180,180,179,179,179,179,180,180,180,180,180,181,181,180,180,181,182,183,183,183,183,182,183,183,183,183,183,183,183,184,185,184,183,183,183,184,184,184,185,185,186,186,185,185,185,186,186,185,184,185,186,185,184,183,183,183,183,182,182,183,184,185,184,183,183,183,184,184,184,184,184,184,185,186,185,184,185,185,185,185,185,184,184,184,184,184,183,183,184,184,184,184,184,185,185,185,184,184,185,185,185,184,184,183,183,183,183,182,182,181,181,181,181,180,180,180,179,179,180,181,181,181,180,180,180,179,178,178,177,176,176,176,176,177,177,177,177,177,176,177,177,176,174,172,173,173,173,172,173,173,173,173,173,173,174,174,174,173,173,173,173,172,171,170,169,168,168,168,168,168,168,168,168,168,168,168,168,
2,2,2,1,2,4,11,17,17,13,10,12,23,36,44,47,52,60,66,66,56,42,32,33,47,75,110,140,157,165,167,168,171,175,176,176,176,175,174,175,176,176,176,176,177,177,175,166,139,94,55,43,48,61,91,133,163,174,175,176,177,177,176,175,176,176,176,177,176,176,176,177,176,177,177,178,179,179,179,178,178,178,178,179,179,179,179,178,178,179,180,180,179,178,180,181,181,181,181,181,181,182,182,182,182,181,181,182,183,184,183,181,180,181,182,182,182,182,182,182,182,181,181,182,182,182,182,181,182,182,182,181,180,181,181,180,179,180,181,182,181,181,181,181,182,182,183,182,181,180,181,182,182,181,181,181,182,182,182,182,181,180,180,181,181,180,180,181,181,181,180,180,180,181,182,182,181,181,181,181,181,181,180,179,179,179,179,179,178,178,178,178,178,178,178,177,177,178,179,179,178,177,177,177,176,176,176,176,175,174,173,173,173,174,174,175,174,173,173,174,173,171,170,170,171,170,170,170,169,169,169,170,171,172,171,171,170,169,169,169,169,168,167,166,165,164,163,164,165,165,165,165,165,165,165,165,
1,1,1,1,2,4,8,12,12,9,8,15,30,46,57,66,68,62,59,60,55,42,31,33,47,70,98,119,130,135,139,146,157,166,170,172,173,172,170,170,172,174,174,174,173,173,171,159,127,79,42,29,30,43,82,133,164,172,173,174,175,175,174,174,175,175,175,175,174,174,175,174,174,174,175,176,177,178,178,177,176,177,177,178,178,178,177,177,177,177,178,177,177,177,179,179,178,177,177,178,179,179,180,180,180,180,180,180,181,182,181,179,178,178,179,179,179,179,179,179,179,179,180,180,180,179,179,179,179,179,179,179,179,179,179,178,178,179,179,179,179,179,179,179,179,180,180,179,179,179,179,180,180,178,178,178,179,179,179,178,178,177,176,176,177,177,178,178,177,177,176,175,176,177,179,180,180,179,178,177,178,177,176,176,176,176,177,177,176,175,175,175,175,175,175,174,173,174,175,175,175,174,174,174,173,174,174,174,174,172,170,169,169,169,170,171,171,171,171,171,170,169,168,169,169,169,168,168,168,167,166,166,168,169,169,168,167,166,165,165,165,165,165,164,164,163,161,162,164,165,165,164,163,163,162,162,
1,1,1,1,2,3,5,6,6,4,6,14,28,41,54,68,70,55,42,41,41,33,29,36,49,66,79,83,86,91,99,115,134,151,160,164,165,162,158,157,163,170,172,171,171,171,169,155,118,67,30,18,21,39,83,134,162,170,171,173,174,174,173,173,174,173,173,173,173,173,173,173,172,172,173,174,175,177,177,176,175,175,176,177,177,177,177,176,175,175,175,175,175,176,178,178,176,174,175,175,176,177,177,178,177,177,177,178,178,179,179,177,176,176,176,176,176,176,176,176,177,177,178,178,178,178,178,177,177,177,177,178,178,178,177,176,177,178,177,176,176,177,177,176,176,176,175,175,177,178,178,178,177,176,175,175,176,177,176,175,174,174,173,174,174,175,177,176,175,174,173,172,172,174,176,178,178,177,176,175,175,175,174,174,174,175,175,175,174,174,174,173,173,173,173,172,171,172,173,174,173,173,172,172,171,172,173,173,173,171,169,167,167,168,168,169,170,170,169,169,168,168,168,168,169,168,168,168,168,167,165,165,165,166,167,166,165,164,163,163,163,164,164,164,163,163,162,162,163,165,165,163,162,161,160,161,
1,1,1,1,2,2,3,3,3,2,4,11,19,26,36,49,52,41,27,23,24,21,22,31,43,53,54,50,51,59,72,88,110,133,146,148,146,139,134,139,153,164,169,170,169,169,166,150,110,57,22,13,20,47,96,140,162,168,171,172,173,173,172,172,172,172,172,172,172,172,172,171,171,172,172,173,174,175,175,174,174,174,174,175,175,175,175,175,173,173,173,174,174,175,177,177,176,175,175,175,175,176,176,176,175,175,175,176,177,178,176,175,174,174,174,174,174,174,174,175,176,176,177,177,177,177,176,175,174,175,176,176,176,176,175,175,175,176,175,173,173,175,175,174,174,173,172,173,175,176,177,176,175,174,174,174,175,175,174,173,172,171,172,173,173,175,177,176,175,173,172,171,170,171,173,175,175,175,174,174,174,174,173,174,174,174,174,174,173,173,173,173,172,172,172,172,171,172,173,174,173,172,172,171,171,171,172,172,171,170,169,168,168,168,168,169,169,170,169,168,167,168,168,168,167,167,167,168,168,167,166,164,164,164,165,165,164,164,163,163,163,163,164,164,164,163,162,162,162,163,163,162,161,159,159,160,
1,1,1,1,1,1,1,1,1,1,3,7,11,14,19,27,31,26,17,14,14,13,15,20,27,33,32,28,33,44,55,67,87,111,121,118,111,103,104,121,144,160,167,168,168,168,164,147,104,51,19,12,23,56,106,146,163,169,171,172,172,172,171,171,171,172,172,172,172,172,171,171,171,171,171,172,172,172,172,172,172,171,172,172,172,173,172,172,171,171,172,173,173,173,175,176,176,175,175,176,176,176,176,175,174,173,173,175,176,176,175,174,173,173,174,174,174,173,173,174,175,176,176,176,176,176,175,174,174,174,175,175,175,175,174,173,173,174,174,172,172,173,173,173,173,172,172,173,175,175,175,174,175,175,174,174,174,174,173,173,171,170,172,173,173,174,176,175,174,173,173,172,170,169,170,171,171,172,172,172,172,172,172,173,174,174,174,173,173,173,173,173,172,172,172,171,171,171,172,173,173,173,172,172,171,171,171,170,169,168,168,168,168,168,168,169,169,170,170,168,168,168,168,167,166,166,167,167,168,167,166,165,163,162,163,163,163,163,163,164,164,163,163,163,163,163,163,162,161,161,162,161,160,160,159,159,
1,1,1,1,1,1,1,1,1,1,2,5,7,9,11,15,18,17,14,12,12,12,11,12,14,17,17,17,22,31,38,47,65,83,87,81,72,65,76,105,135,154,164,167,167,167,165,147,103,51,20,15,30,66,112,147,163,169,171,172,172,171,170,170,172,173,172,172,171,171,171,170,170,170,171,171,170,170,170,170,170,170,170,170,170,171,170,170,169,169,169,170,170,170,171,173,174,175,175,176,176,177,177,176,173,172,173,174,175,175,175,174,174,174,174,174,174,173,173,175,176,177,176,176,176,175,175,175,175,175,175,175,175,175,174,173,173,174,174,173,172,172,172,173,173,173,173,174,175,174,173,173,174,175,174,173,173,173,172,172,171,171,172,172,172,173,174,174,173,173,173,173,172,171,170,170,169,169,170,171,171,171,171,172,173,175,174,173,173,173,173,172,172,172,171,171,171,171,171,171,172,172,172,172,171,171,170,168,168,167,167,167,167,167,167,168,169,169,169,169,168,168,167,166,165,165,165,166,167,167,166,165,163,162,162,162,163,163,163,163,163,162,162,162,162,163,163,162,161,161,161,161,162,161,160,159,
1,1,1,2,2,1,1,1,1,1,2,4,5,6,8,10,13,14,13,12,12,12,11,10,9,10,10,11,15,21,25,31,44,54,55,50,41,37,54,87,118,141,155,161,162,163,165,151,109,56,24,20,40,79,122,151,165,170,172,172,171,171,170,171,172,172,171,170,170,169,168,169,169,169,170,170,170,169,169,170,170,170,170,169,170,170,169,169,169,168,168,168,166,165,166,168,171,173,175,175,176,177,177,175,171,169,171,173,174,175,176,177,176,174,173,174,173,173,173,175,177,178,177,177,176,176,177,177,177,177,176,176,175,175,174,174,174,175,175,174,173,172,173,174,174,174,174,175,174,173,172,172,173,174,174,174,173,171,170,171,172,171,171,171,171,172,172,173,173,173,172,173,173,172,172,171,170,169,170,170,170,169,168,169,172,174,174,173,173,173,173,172,171,171,170,170,171,171,170,170,171,172,172,171,170,170,169,167,167,167,167,167,167,165,166,168,168,168,168,169,168,167,167,166,164,163,163,165,166,166,165,164,163,162,162,163,163,163,163,163,162,162,161,161,162,162,163,162,162,161,161,162,163,163,161,161,
1,1,2,2,2,1,1,1,2,2,2,3,4,5,6,8,10,12,12,11,10,11,10,9,8,8,9,10,12,15,18,24,31,33,30,27,22,22,37,64,93,118,135,142,143,147,156,152,117,62,27,27,52,94,134,158,167,170,171,171,171,170,170,171,171,171,171,170,169,168,166,167,168,168,169,170,170,169,169,170,171,171,170,170,170,170,169,169,169,169,169,168,166,164,163,165,170,173,175,176,177,177,176,174,169,167,169,173,174,175,177,178,177,174,173,173,173,172,172,174,177,179,179,179,180,180,180,181,181,180,178,176,174,174,175,176,176,175,174,173,173,173,174,174,175,175,174,174,174,173,172,172,173,174,174,175,174,171,169,170,172,172,171,171,172,173,173,174,174,173,172,173,173,172,172,171,171,170,170,169,169,169,168,168,170,172,172,172,173,173,173,172,171,170,170,170,171,172,172,172,172,173,172,170,169,169,169,168,168,168,168,168,167,165,166,167,168,168,168,168,168,168,167,166,165,165,164,165,166,166,165,164,164,164,165,165,165,165,165,164,163,163,163,163,163,163,163,163,163,163,163,164,165,165,164,163,
1,2,2,2,2,2,2,2,3,3,3,4,5,5,6,7,9,10,10,9,10,10,9,7,7,9,11,11,12,13,15,22,26,22,15,12,12,15,27,47,71,94,107,108,109,120,137,142,114,63,30,35,69,111,145,163,168,170,170,170,170,170,170,170,171,172,172,171,171,169,169,169,169,169,170,171,170,170,170,171,172,172,171,171,171,170,169,169,171,172,171,171,170,168,167,168,171,174,177,177,177,176,175,174,171,169,171,174,175,175,176,177,176,173,173,175,174,172,171,173,176,179,181,182,183,184,184,184,184,183,180,176,174,174,175,176,177,176,174,174,174,174,175,175,176,175,174,174,175,175,174,173,173,174,174,175,175,173,170,170,172,173,173,173,174,175,176,176,175,174,174,174,173,173,172,173,172,172,171,170,170,170,170,171,172,173,173,173,173,173,173,172,172,173,173,172,172,173,174,175,176,175,174,172,171,171,171,170,170,169,169,169,168,168,168,169,169,169,168,168,168,168,169,169,168,168,168,168,169,168,168,167,168,168,167,168,168,168,167,166,165,166,167,167,166,165,164,164,164,165,164,165,166,166,166,166,
1,1,2,2,3,4,5,4,4,4,4,5,5,6,6,7,8,8,8,10,13,13,10,7,7,10,14,15,14,13,15,19,20,14,7,6,9,13,22,36,54,72,78,73,77,96,115,117,94,57,36,52,94,134,158,167,169,170,170,170,170,170,171,171,172,173,174,173,173,172,172,172,172,171,171,171,171,172,173,174,174,173,173,173,172,170,170,171,173,174,173,173,173,173,173,173,174,176,177,178,178,178,177,176,175,174,175,176,177,177,177,177,176,175,175,176,176,174,174,175,176,178,180,182,183,185,185,185,185,183,180,177,175,175,176,176,177,177,176,176,177,177,177,177,177,176,176,176,176,177,176,176,175,175,175,177,177,175,173,172,174,175,176,175,176,178,178,178,177,176,176,176,175,174,175,176,175,175,175,174,174,174,174,175,176,177,176,175,175,175,174,174,175,176,176,175,174,174,176,177,178,178,177,176,174,174,174,173,172,172,171,171,171,171,171,170,170,171,171,170,170,170,170,171,171,171,171,171,172,172,171,171,171,170,170,170,170,170,169,167,167,167,169,169,169,167,166,165,165,166,166,165,166,167,168,168,
1,1,2,2,4,6,8,8,6,5,5,6,6,7,7,8,8,8,9,12,16,15,10,6,7,12,17,19,17,15,15,16,13,8,5,6,9,12,18,25,35,48,54,52,60,84,99,90,66,45,45,76,122,155,168,170,171,171,172,172,172,172,172,172,173,174,175,175,174,173,174,174,174,172,171,172,172,173,175,176,176,175,174,174,174,172,171,173,175,175,174,174,175,176,176,176,176,176,177,178,179,179,179,178,177,177,177,178,179,179,178,178,178,177,178,178,178,177,177,177,177,178,180,180,181,182,182,183,182,181,180,179,178,178,178,178,178,178,179,179,179,179,179,179,179,179,178,178,178,178,178,179,179,178,178,178,178,177,175,175,176,178,178,177,178,179,179,179,178,178,178,177,176,176,177,178,178,178,179,178,178,178,178,179,179,179,178,177,177,177,176,176,178,179,179,177,176,175,176,177,178,178,178,177,176,176,176,175,174,173,173,173,173,173,172,171,172,173,173,172,171,171,171,172,173,173,172,172,172,173,173,173,172,171,171,171,171,170,169,168,168,168,168,169,169,169,167,166,166,166,166,166,166,167,168,168,
1,1,2,2,4,6,9,10,8,6,6,6,6,7,8,8,8,8,9,13,17,15,9,6,7,13,19,21,18,15,15,14,10,5,4,6,9,12,15,19,25,36,43,45,56,81,94,79,52,38,50,90,136,164,171,171,171,172,173,173,174,174,173,172,173,175,176,176,174,173,174,175,174,173,172,172,173,174,176,177,176,175,175,175,175,173,172,174,176,175,174,175,175,176,177,177,177,176,176,178,179,180,180,179,178,178,178,179,180,180,179,179,179,179,179,179,178,178,179,178,178,179,180,180,179,180,181,181,181,180,180,179,180,180,179,178,178,179,180,180,180,180,181,180,180,180,179,179,178,178,179,181,181,180,179,179,178,177,176,176,177,178,179,178,178,179,180,179,178,178,178,178,176,176,178,179,179,179,180,180,180,179,179,180,180,180,179,178,178,178,177,177,179,180,179,177,176,176,176,177,178,178,178,177,176,176,177,176,175,174,174,173,173,173,172,172,172,174,174,173,171,171,172,173,173,173,172,172,171,172,173,173,172,171,171,171,171,170,169,169,168,167,167,168,169,169,168,167,166,166,166,166,166,167,168,168
);
signal counter : integer range 0 to 1000;
signal c : integer range 0 to 65535 :=0;
signal d : integer range 0 to 65535 :=0;
signal test: integer range 0 to 255:=0;
signal testdata: std_logic_vector(7 downto 0):="00000000";
signal Xpos,Ypos: integer range 0 to 799:=0;
---------------------------sync-----------------------------
signal BUFF_WAIT: std_logic:='0';
signal VGAFLAG: std_logic_vector(2 downto 0);
-------------------------ram/gray----------------------------
signal RAMFULL_POINTER:integer range 0 to 511:=0;
signal RAMRESTART_POINTER: integer range 0 to 511:=0;
signal RAMADDR1GR,RAMADDR2GR: std_logic_vector(8 downto 0):=(others=>'0');
signal RAMADDR1GR_sync0,RAMADDR1GR_sync1,RAMADDR1GR_sync2,RAMADDR1_bin: std_logic_vector(8 downto 0);
signal RAMADDR2GR_sync0,RAMADDR2GR_sync1,RAMADDR2GR_sync2,RAMADDR2_bin: std_logic_vector(8 downto 0);
-------------------------dual ram ----------------------------------
signal RAMIN1,RAMIN2,RAMOUT1,RAMOUT2: std_logic_vector(7 downto 0);
signal RAMWE1,RAMWE2: std_logic:='0';
signal RAMADDR1,RAMADDR2: integer range 0 to 511:=0;
------------------vga----------------------------------
signal NEXTFRAME: std_logic_vector(2 downto 0):="000";
signal FRAMEEND,FRAMESTART: std_logic:='0';
signal ACTVIDEO: std_logic:='0';
signal VGABEGIN: std_logic:='0';
signal RED,GREEN,BLUE: STD_LOGIC_VECTOR(7 downto 0);
------------------clock--------------------------------
SIGNAL CLK143,CLK143_2,CLK49_5: STD_LOGIC;
------------------sdram--------------------------------
SIGNAL SDRAM_ADDR: STD_LOGIC_VECTOR(24 downto 0);
SIGNAL SDRAM_BE_N: STD_LOGIC_VECTOR(1 downto 0);
SIGNAL SDRAM_CS: STD_LOGIC;
SIGNAL SDRAM_RDVAL,SDRAM_WAIT:STD_LOGIC;
SIGNAL SDRAM_RE_N,SDRAM_WE_N: STD_LOGIC;
SIGNAL SDRAM_READDATA,SDRAM_WRITEDATA: STD_LOGIC_VECTOR(15 downto 0);
SIGNAL DRAM_DQM : STD_LOGIC_VECTOR(1 downto 0);

--------------------------------------------------------

	component true_dual_port_ram_dual_clock is
	port 
	(
		clk_a	: in std_logic;
		clk_b	: in std_logic;
		addr_a	: in natural range 0 to 511;
		addr_b	: in natural range 0 to 511;
		data_a	: in std_logic_vector(7 downto 0);
		data_b	: in std_logic_vector(7 downto 0);
		we_a	: in std_logic := '1';
		we_b	: in std_logic := '1';
		q_a		: out std_logic_vector(7 downto 0);
		q_b		: out std_logic_vector(7 downto 0)
	);
	end component true_dual_port_ram_dual_clock;
   component  vga is
	port(
		CLK: in std_logic;
		R_OUT,G_OUT,B_OUT: OUT std_logic_vector(7 downto 0);
		R_IN,G_IN,B_IN: IN std_logic_vector(7 downto 0);
		VGAHS, VGAVS:OUT std_logic;
	   ACTVID: OUT std_logic;
		VGA_FRAMESTART: out std_logic;
		VGA_FRAMEEND: out std_logic
	);
end component vga;


component ramsys is
        port (
            clk_clk             : in    std_logic                     := 'X';             -- clk
            reset_reset_n       : in    std_logic                     := 'X';             -- reset_n
            clk143_shift_clk    : out   std_logic;                                        -- clk
            clk143_clk          : out   std_logic;                                        -- clk
            clk49_5_clk         : out   std_logic;                                        -- clk
            wire_addr           : out   std_logic_vector(12 downto 0);                    -- addr
            wire_ba             : out   std_logic_vector(1 downto 0);                     -- ba
            wire_cas_n          : out   std_logic;                                        -- cas_n
            wire_cke            : out   std_logic;                                        -- cke
            wire_cs_n           : out   std_logic;                                        -- cs_n
            wire_dq             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
            wire_dqm            : out   std_logic_vector(1 downto 0);                     -- dqm
            wire_ras_n          : out   std_logic;                                        -- ras_n
            wire_we_n           : out   std_logic;                                        -- we_n
            sdram_address       : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
            sdram_byteenable_n  : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
            sdram_chipselect    : in    std_logic                     := 'X';             -- chipselect
            sdram_writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
            sdram_read_n        : in    std_logic                     := 'X';             -- read_n
            sdram_write_n       : in    std_logic                     := 'X';             -- write_n
            sdram_readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
            sdram_readdatavalid : out   std_logic;                                        -- readdatavalid
            sdram_waitrequest   : out   std_logic                                         -- waitrequest
        );
    end component ramsys;
begin


	u0 : component ramsys
        port map (
            clk_clk             => CLOCK_50,             --          clk.clk
            reset_reset_n       => '1',       --        reset.reset_n
            clk143_shift_clk    => CLK143_2,    -- clk143_shift.clk
            clk143_clk          => CLK143,          --       clk143.clk
            clk49_5_clk         => CLK49_5,         --      clk49_5.clk
            wire_addr           => DRAM_ADDR,           --         wire.addr
            wire_ba             => DRAM_BA,             --             .ba
            wire_cas_n          => DRAM_CAS_N,          --             .cas_n
            wire_cke            => DRAM_CKE,            --             .cke
            wire_cs_n           => DRAM_CS_N,           --             .cs_n
            wire_dq             => DRAM_DQ,             --             .dq
            wire_dqm            => DRAM_DQM,            --             .dqm
            wire_ras_n          => DRAM_RAS_N,          --             .ras_n
            wire_we_n           => DRAM_WE_N,           --             .we_n
            sdram_address       => SDRAM_ADDR,       --        sdram.address
            sdram_byteenable_n  => SDRAM_BE_N,  --             .byteenable_n
            sdram_chipselect    => SDRAM_CS,    --             .chipselect
            sdram_writedata     => SDRAM_WRITEDATA,     --             .writedata
            sdram_read_n        => SDRAM_RE_N,        --             .read_n
            sdram_write_n       => SDRAM_WE_N,       --             .write_n
            sdram_readdata      => SDRAM_READDATA,      --             .readdata
            sdram_readdatavalid => SDRAM_RDVAL, --             .readdatavalid
            sdram_waitrequest   => SDRAM_WAIT    --             .waitrequest
        );

      u1 : component vga 
			port map(
					CLK=>CLK49_5,
					R_OUT=>VGA_R,
					G_OUT=>VGA_G,
					B_OUT=>VGA_B,
					R_IN=>RED,
					G_IN=>GREEN,
					B_IN=>BLUE,
					VGAHS=>VGA_HS,
					VGAVS=>VGA_VS,
				   ACTVID=>ACTVIDEO,
					VGA_FRAMESTART=>FRAMESTART,
					VGA_FRAMEEND=>FRAMEEND
			);

		u3: component true_dual_port_ram_dual_clock
		   port map  (
			clk_a=>CLK143,
			clk_b=>clk49_5,
			addr_a=>RAMADDR1,
			addr_b=>RAMADDR2,
			data_a=>RAMIN1,
			data_b=>RAMIN2,
			we_a=>RAMWE1,
			we_b=>RAMWE2,
			q_a=>RAMOUT1,
			q_b=>RAMOUT2			
			);





DRAM_LDQM<=DRAM_DQM(0);
DRAM_UDQM<=DRAM_DQM(1);
DRAM_CLK<=CLK143_2;
VGA_CLK<=CLK49_5;
SDRAM_CS<='1';
SDRAM_BE_N<="00";
VGA_BLANK_N<='1';
VGA_SYNC_N<='0';
ilk: PROCESS (CLK143)
begin
if rising_edge(clk143)then
------------double flop sync----------------------
	RAMADDR2GR_sync0<=RAMADDR2GR;
	RAMADDR2GR_sync1<=RAMADDR2GR_sync0;
	RAMADDR2_bin<=gray_to_bin(RAMADDR2GR_sync1);
   NEXTFRAME(1)<=NEXTFRAME(0);
	NEXTFRAME(2)<=NEXTFRAME(1);


RAMADDR1GR<=bin_to_gray(std_logic_vector(to_unsigned(RAMADDR1,9)));
----------------------------------------------------
	case BUFF_CTRL is
		when st0=>------------write image to  SDRAM     
		if (SDRAM_WAIT='0')then	
		    SDRAM_WE_N<='0';
			 SDRAM_RE_N<='1';
------------------------circle generation------------------
				if(Xpos<799)then
					Xpos<=Xpos+1;
				else
					Xpos<=0;
				  if(Ypos<599)then
						Ypos<=Ypos+1;
				  else
						Ypos<=0;
				  end if;	  
				end if;
				IF((Xpos > 10 and Xpos < 267) and(Ypos > 200 and Ypos < 457) )THEN
					test<=Rom(c);
					c <= c + 1;
				elsif((Xpos > 280 and Xpos < 537) and(Ypos > 200 and Ypos < 457) )THEN
					test<=ROM_Gauss(d);
					d <= d + 1;
				else
					test<=0;
				end if;
				
			
				
------------------------------------------------------------
			 SDRAM_WRITEDATA(7 downto 0) <= std_logic_vector(to_unsigned(test, 8));
	       SDRAM_ADDR<=std_logic_vector(unsigned(SDRAM_ADDR)+1);	

		end if;	
		
      if(to_integer(unsigned(SDRAM_ADDR))>(800*600-1) )then-----800x600 resolution
		   RAMADDR1<=0;
			BUFF_WAIT<='0';
			RAMFULL_POINTER<=10;----------min. value 2
		   BUFF_CTRL<=st1;
			SDRAM_ADDR<=(others=>'0');
		end if;
		
		when st1=>-----------write from SDRAM to BUFFER
		      SDRAM_WE_N<='1';
            RAMWE1<=SDRAM_RDVAL;
			IF(BUFF_WAIT='0')then
					 SDRAM_RE_N<='0';
					   ------------if no wait request is issued and read enable------
		            IF(SDRAM_WAIT='0' and SDRAM_RE_N='0')THEN	
							IF(RAMFULL_POINTER<511)then-----move full pointer
								RAMFULL_POINTER<=RAMFULL_POINTER+1;
								else
								RAMFULL_POINTER<=0;
							end if;			
			            SDRAM_ADDR<=std_logic_vector(unsigned(SDRAM_ADDR)+1);		
	               END IF;
						-------------check if the buffer is full----------------------
						IF(to_integer(unsigned(RAMADDR2_bin))=(RAMFULL_POINTER))then
								VGAFLAG(0)<='1';---------init displaying image
								SDRAM_RE_N<='1';
								BUFF_WAIT<='1';
								IF((RAMADDR2+63)<511)THEN
									RAMRESTART_POINTER<=to_integer(unsigned(RAMADDR2_bin))+63;
									ELSE
									RAMRESTART_POINTER<=to_integer(unsigned(RAMADDR2_bin))+63-511;
								END IF;
						end if;
			END IF;
			    	RAMIN1<=SDRAM_READDATA(7 downto 0);	
					------------while data is avalable, write to buffer RAM
					IF(SDRAM_RDVAL='1')then
						IF(RAMADDR1<511)then
						RAMADDR1<=RAMADDR1+1;
						else
						RAMADDR1<=0;
						end if;
					END IF;
					-------------------------------refill buffer------------------------
					     IF(to_integer(unsigned(RAMADDR2_bin))=RAMRESTART_POINTER and BUFF_WAIT='1')then
						  BUFF_WAIT<='0';		  
						  end if;
					-------------------------------end of frame--------------------------
 				        IF(NEXTFRAME(2)='1')THEN
						      xpos<=0;
	                    	ypos<=0;
							   BUFF_CTRL<=ST0;
								VGAFLAG(0)<='0';
								SDRAM_ADDR<=(others=>'0');
								------------
								counter<=0;
								test<=0;
							END IF;
		    
		when others=>NULL;
		END CASE;





end if;
end process ilk;
ilk_i: PROCESS(CLK49_5)
begin
if rising_edge(CLK49_5)then
	 
RAMADDR2GR<=bin_to_gray(std_logic_vector(to_unsigned(RAMADDR2,9)));
-------------dual clock sync-------------------------
RAMADDR1GR_sync0<=RAMADDR1GR;
RAMADDR1GR_sync1<=RAMADDR1GR_sync0;
VGAFLAG(1)<=VGAFLAG(0);
VGAFLAG(2)<=VGAFLAG(1);

RAMADDR1_bin<=gray_to_bin(RAMADDR1GR_sync1);


    IF(VGAFLAG(2)='1' AND FRAMESTART='1' )THEN-------if buffer is rdy and  begin of new frame, start displaying image
	 VGABEGIN<='1';
	 end if;
	 
	 IF(FRAMEEND='1' AND VGABEGIN='1')THEN------end of frame
	 NEXTFRAME(0)<='1';
	 VGABEGIN<='0';
	 ELSE
	 NEXTFRAME(0)<='0';
	 END IF;
	
		IF(ACTVIDEO='1'AND to_integer(unsigned(RAMADDR1_bin))/=RAMADDR2  AND VGABEGIN='1')then----if buffer ia not empty
			IF(RAMADDR2<511)then
			RAMADDR2<=RAMADDR2+1;
			else
			RAMADDR2<=0;
			end if;
		   RED<=RAMOUT2;
	      GREEN<=RAMOUT2;
		   BLUE<=RAMOUT2;
		ELSIF(VGABEGIN='0')THEN---------if buffer not ready
	   RAMADDR2<=0;
		BLUE<=(others=>'0');
		RED<=(others=>'0');
		GREEN<=(others=>'0');
		END IF;
end if;
end process ilk_i ;
-----------------------------------------------------------------------------------

-----------------------------------------------------------------------------------
end main;